module mime

fn load_data() map[string]MimeType {
    mut data := map[string]MimeType{}
    data['application/1d-interleaved-parityfec'] = MimeType{'iana',[]string,false,''}
    data['application/3gpdash-qoe-report+xml'] = MimeType{'iana',[]string,true,''}
    data['application/3gpp-ims+xml'] = MimeType{'iana',[]string,true,''}
    data['application/a2l'] = MimeType{'iana',[]string,false,''}
    data['application/activemessage'] = MimeType{'iana',[]string,false,''}
    data['application/activity+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-costmap+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-costmapfilter+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-directory+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-endpointcost+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-endpointcostparams+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-endpointprop+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-endpointpropparams+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-error+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-networkmap+json'] = MimeType{'iana',[]string,true,''}
    data['application/alto-networkmapfilter+json'] = MimeType{'iana',[]string,true,''}
    data['application/aml'] = MimeType{'iana',[]string,false,''}
    data['application/andrew-inset'] = MimeType{'iana',['ez'],false,''}
    data['application/applefile'] = MimeType{'iana',[]string,false,''}
    data['application/applixware'] = MimeType{'apache',['aw'],false,''}
    data['application/atf'] = MimeType{'iana',[]string,false,''}
    data['application/atfx'] = MimeType{'iana',[]string,false,''}
    data['application/atom+xml'] = MimeType{'iana',['atom'],true,''}
    data['application/atomcat+xml'] = MimeType{'iana',['atomcat'],true,''}
    data['application/atomdeleted+xml'] = MimeType{'iana',[]string,true,''}
    data['application/atomicmail'] = MimeType{'iana',[]string,false,''}
    data['application/atomsvc+xml'] = MimeType{'iana',['atomsvc'],true,''}
    data['application/atsc-dwd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/atsc-held+xml'] = MimeType{'iana',[]string,true,''}
    data['application/atsc-rsat+xml'] = MimeType{'iana',[]string,true,''}
    data['application/atxml'] = MimeType{'iana',[]string,false,''}
    data['application/auth-policy+xml'] = MimeType{'iana',[]string,true,''}
    data['application/bacnet-xdd+zip'] = MimeType{'iana',[]string,false,''}
    data['application/batch-smtp'] = MimeType{'iana',[]string,false,''}
    data['application/bdoc'] = MimeType{'',['bdoc'],false,''}
    data['application/beep+xml'] = MimeType{'iana',[]string,true,''}
    data['application/calendar+json'] = MimeType{'iana',[]string,true,''}
    data['application/calendar+xml'] = MimeType{'iana',[]string,true,''}
    data['application/call-completion'] = MimeType{'iana',[]string,false,''}
    data['application/cals-1840'] = MimeType{'iana',[]string,false,''}
    data['application/cbor'] = MimeType{'iana',[]string,false,''}
    data['application/cccex'] = MimeType{'iana',[]string,false,''}
    data['application/ccmp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/ccxml+xml'] = MimeType{'iana',['ccxml'],true,''}
    data['application/cdfx+xml'] = MimeType{'iana',[]string,true,''}
    data['application/cdmi-capability'] = MimeType{'iana',['cdmia'],false,''}
    data['application/cdmi-container'] = MimeType{'iana',['cdmic'],false,''}
    data['application/cdmi-domain'] = MimeType{'iana',['cdmid'],false,''}
    data['application/cdmi-object'] = MimeType{'iana',['cdmio'],false,''}
    data['application/cdmi-queue'] = MimeType{'iana',['cdmiq'],false,''}
    data['application/cdni'] = MimeType{'iana',[]string,false,''}
    data['application/cea'] = MimeType{'iana',[]string,false,''}
    data['application/cea-2018+xml'] = MimeType{'iana',[]string,true,''}
    data['application/cellml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/cfw'] = MimeType{'iana',[]string,false,''}
    data['application/clue_info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/cms'] = MimeType{'iana',[]string,false,''}
    data['application/cnrp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/coap-group+json'] = MimeType{'iana',[]string,true,''}
    data['application/coap-payload'] = MimeType{'iana',[]string,false,''}
    data['application/commonground'] = MimeType{'iana',[]string,false,''}
    data['application/conference-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/cose'] = MimeType{'iana',[]string,false,''}
    data['application/cose-key'] = MimeType{'iana',[]string,false,''}
    data['application/cose-key-set'] = MimeType{'iana',[]string,false,''}
    data['application/cpl+xml'] = MimeType{'iana',[]string,true,''}
    data['application/csrattrs'] = MimeType{'iana',[]string,false,''}
    data['application/csta+xml'] = MimeType{'iana',[]string,true,''}
    data['application/cstadata+xml'] = MimeType{'iana',[]string,true,''}
    data['application/csvm+json'] = MimeType{'iana',[]string,true,''}
    data['application/cu-seeme'] = MimeType{'apache',['cu'],false,''}
    data['application/cwt'] = MimeType{'iana',[]string,false,''}
    data['application/cybercash'] = MimeType{'iana',[]string,false,''}
    data['application/dart'] = MimeType{'',[]string,true,''}
    data['application/dash+xml'] = MimeType{'iana',['mpd'],true,''}
    data['application/dashdelta'] = MimeType{'iana',[]string,false,''}
    data['application/davmount+xml'] = MimeType{'iana',['davmount'],true,''}
    data['application/dca-rft'] = MimeType{'iana',[]string,false,''}
    data['application/dcd'] = MimeType{'iana',[]string,false,''}
    data['application/dec-dx'] = MimeType{'iana',[]string,false,''}
    data['application/dialog-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/dicom'] = MimeType{'iana',[]string,false,''}
    data['application/dicom+json'] = MimeType{'iana',[]string,true,''}
    data['application/dicom+xml'] = MimeType{'iana',[]string,true,''}
    data['application/dii'] = MimeType{'iana',[]string,false,''}
    data['application/dit'] = MimeType{'iana',[]string,false,''}
    data['application/dns'] = MimeType{'iana',[]string,false,''}
    data['application/dns+json'] = MimeType{'iana',[]string,true,''}
    data['application/dns-message'] = MimeType{'iana',[]string,false,''}
    data['application/docbook+xml'] = MimeType{'apache',['dbk'],true,''}
    data['application/dskpp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/dssc+der'] = MimeType{'iana',['dssc'],false,''}
    data['application/dssc+xml'] = MimeType{'iana',['xdssc'],true,''}
    data['application/dvcs'] = MimeType{'iana',[]string,false,''}
    data['application/ecmascript'] = MimeType{'iana',['ecma', 'es'],true,''}
    data['application/edi-consent'] = MimeType{'iana',[]string,false,''}
    data['application/edi-x12'] = MimeType{'iana',[]string,false,''}
    data['application/edifact'] = MimeType{'iana',[]string,false,''}
    data['application/efi'] = MimeType{'iana',[]string,false,''}
    data['application/emergencycalldata.comment+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emergencycalldata.control+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emergencycalldata.deviceinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emergencycalldata.ecall.msd'] = MimeType{'iana',[]string,false,''}
    data['application/emergencycalldata.providerinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emergencycalldata.serviceinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emergencycalldata.subscriberinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emergencycalldata.veds+xml'] = MimeType{'iana',[]string,true,''}
    data['application/emma+xml'] = MimeType{'iana',['emma'],true,''}
    data['application/emotionml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/encaprtp'] = MimeType{'iana',[]string,false,''}
    data['application/epp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/epub+zip'] = MimeType{'iana',['epub'],false,''}
    data['application/eshop'] = MimeType{'iana',[]string,false,''}
    data['application/exi'] = MimeType{'iana',['exi'],false,''}
    data['application/expect-ct-report+json'] = MimeType{'iana',[]string,true,''}
    data['application/fastinfoset'] = MimeType{'iana',[]string,false,''}
    data['application/fastsoap'] = MimeType{'iana',[]string,false,''}
    data['application/fdt+xml'] = MimeType{'iana',[]string,true,''}
    data['application/fhir+json'] = MimeType{'iana',[]string,true,''}
    data['application/fhir+xml'] = MimeType{'iana',[]string,true,''}
    data['application/fido.trusted-apps+json'] = MimeType{'',[]string,true,''}
    data['application/fits'] = MimeType{'iana',[]string,false,''}
    data['application/font-sfnt'] = MimeType{'iana',[]string,false,''}
    data['application/font-tdpfr'] = MimeType{'iana',['pfr'],false,''}
    data['application/font-woff'] = MimeType{'iana',[]string,false,''}
    data['application/framework-attributes+xml'] = MimeType{'iana',[]string,true,''}
    data['application/geo+json'] = MimeType{'iana',['geojson'],true,''}
    data['application/geo+json-seq'] = MimeType{'iana',[]string,false,''}
    data['application/geopackage+sqlite3'] = MimeType{'iana',[]string,false,''}
    data['application/geoxacml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/gltf-buffer'] = MimeType{'iana',[]string,false,''}
    data['application/gml+xml'] = MimeType{'iana',['gml'],true,''}
    data['application/gpx+xml'] = MimeType{'apache',['gpx'],true,''}
    data['application/gxf'] = MimeType{'apache',['gxf'],false,''}
    data['application/gzip'] = MimeType{'iana',['gz'],false,''}
    data['application/h224'] = MimeType{'iana',[]string,false,''}
    data['application/held+xml'] = MimeType{'iana',[]string,true,''}
    data['application/hjson'] = MimeType{'',['hjson'],false,''}
    data['application/http'] = MimeType{'iana',[]string,false,''}
    data['application/hyperstudio'] = MimeType{'iana',['stk'],false,''}
    data['application/ibe-key-request+xml'] = MimeType{'iana',[]string,true,''}
    data['application/ibe-pkg-reply+xml'] = MimeType{'iana',[]string,true,''}
    data['application/ibe-pp-data'] = MimeType{'iana',[]string,false,''}
    data['application/iges'] = MimeType{'iana',[]string,false,''}
    data['application/im-iscomposing+xml'] = MimeType{'iana',[]string,true,''}
    data['application/index'] = MimeType{'iana',[]string,false,''}
    data['application/index.cmd'] = MimeType{'iana',[]string,false,''}
    data['application/index.obj'] = MimeType{'iana',[]string,false,''}
    data['application/index.response'] = MimeType{'iana',[]string,false,''}
    data['application/index.vnd'] = MimeType{'iana',[]string,false,''}
    data['application/inkml+xml'] = MimeType{'iana',['ink', 'inkml'],true,''}
    data['application/iotp'] = MimeType{'iana',[]string,false,''}
    data['application/ipfix'] = MimeType{'iana',['ipfix'],false,''}
    data['application/ipp'] = MimeType{'iana',[]string,false,''}
    data['application/isup'] = MimeType{'iana',[]string,false,''}
    data['application/its+xml'] = MimeType{'iana',[]string,true,''}
    data['application/java-archive'] = MimeType{'apache',['jar', 'war', 'ear'],false,''}
    data['application/java-serialized-object'] = MimeType{'apache',['ser'],false,''}
    data['application/java-vm'] = MimeType{'apache',['class'],false,''}
    data['application/javascript'] = MimeType{'iana',['js', 'mjs'],true,'UTF-8'}
    data['application/jf2feed+json'] = MimeType{'iana',[]string,true,''}
    data['application/jose'] = MimeType{'iana',[]string,false,''}
    data['application/jose+json'] = MimeType{'iana',[]string,true,''}
    data['application/jrd+json'] = MimeType{'iana',[]string,true,''}
    data['application/json'] = MimeType{'iana',['json', 'map'],true,'UTF-8'}
    data['application/json-patch+json'] = MimeType{'iana',[]string,true,''}
    data['application/json-seq'] = MimeType{'iana',[]string,false,''}
    data['application/json5'] = MimeType{'',['json5'],false,''}
    data['application/jsonml+json'] = MimeType{'apache',['jsonml'],true,''}
    data['application/jwk+json'] = MimeType{'iana',[]string,true,''}
    data['application/jwk-set+json'] = MimeType{'iana',[]string,true,''}
    data['application/jwt'] = MimeType{'iana',[]string,false,''}
    data['application/kpml-request+xml'] = MimeType{'iana',[]string,true,''}
    data['application/kpml-response+xml'] = MimeType{'iana',[]string,true,''}
    data['application/ld+json'] = MimeType{'iana',['jsonld'],true,''}
    data['application/lgr+xml'] = MimeType{'iana',[]string,true,''}
    data['application/link-format'] = MimeType{'iana',[]string,false,''}
    data['application/load-control+xml'] = MimeType{'iana',[]string,true,''}
    data['application/lost+xml'] = MimeType{'iana',['lostxml'],true,''}
    data['application/lostsync+xml'] = MimeType{'iana',[]string,true,''}
    data['application/lxf'] = MimeType{'iana',[]string,false,''}
    data['application/mac-binhex40'] = MimeType{'iana',['hqx'],false,''}
    data['application/mac-compactpro'] = MimeType{'apache',['cpt'],false,''}
    data['application/macwriteii'] = MimeType{'iana',[]string,false,''}
    data['application/mads+xml'] = MimeType{'iana',['mads'],true,''}
    data['application/manifest+json'] = MimeType{'',['webmanifest'],true,'UTF-8'}
    data['application/marc'] = MimeType{'iana',['mrc'],false,''}
    data['application/marcxml+xml'] = MimeType{'iana',['mrcx'],true,''}
    data['application/mathematica'] = MimeType{'iana',['ma', 'nb', 'mb'],false,''}
    data['application/mathml+xml'] = MimeType{'iana',['mathml'],true,''}
    data['application/mathml-content+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mathml-presentation+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-associated-procedure-description+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-deregister+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-envelope+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-msk+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-msk-response+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-protection-description+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-reception-report+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-register+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-register-response+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-schedule+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbms-user-service-description+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mbox'] = MimeType{'iana',['mbox'],false,''}
    data['application/media-policy-dataset+xml'] = MimeType{'iana',[]string,true,''}
    data['application/media_control+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mediaservercontrol+xml'] = MimeType{'iana',['mscml'],true,''}
    data['application/merge-patch+json'] = MimeType{'iana',[]string,true,''}
    data['application/metalink+xml'] = MimeType{'apache',['metalink'],true,''}
    data['application/metalink4+xml'] = MimeType{'iana',['meta4'],true,''}
    data['application/mets+xml'] = MimeType{'iana',['mets'],true,''}
    data['application/mf4'] = MimeType{'iana',[]string,false,''}
    data['application/mikey'] = MimeType{'iana',[]string,false,''}
    data['application/mmt-aei+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mmt-usd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mods+xml'] = MimeType{'iana',['mods'],true,''}
    data['application/moss-keys'] = MimeType{'iana',[]string,false,''}
    data['application/moss-signature'] = MimeType{'iana',[]string,false,''}
    data['application/mosskey-data'] = MimeType{'iana',[]string,false,''}
    data['application/mosskey-request'] = MimeType{'iana',[]string,false,''}
    data['application/mp21'] = MimeType{'iana',['m21', 'mp21'],false,''}
    data['application/mp4'] = MimeType{'iana',['mp4s', 'm4p'],false,''}
    data['application/mpeg4-generic'] = MimeType{'iana',[]string,false,''}
    data['application/mpeg4-iod'] = MimeType{'iana',[]string,false,''}
    data['application/mpeg4-iod-xmt'] = MimeType{'iana',[]string,false,''}
    data['application/mrb-consumer+xml'] = MimeType{'iana',[]string,true,''}
    data['application/mrb-publish+xml'] = MimeType{'iana',[]string,true,''}
    data['application/msc-ivr+xml'] = MimeType{'iana',[]string,true,''}
    data['application/msc-mixer+xml'] = MimeType{'iana',[]string,true,''}
    data['application/msword'] = MimeType{'iana',['doc', 'dot'],false,''}
    data['application/mud+json'] = MimeType{'iana',[]string,true,''}
    data['application/mxf'] = MimeType{'iana',['mxf'],false,''}
    data['application/n-quads'] = MimeType{'iana',['nq'],false,''}
    data['application/n-triples'] = MimeType{'iana',['nt'],false,''}
    data['application/nasdata'] = MimeType{'iana',[]string,false,''}
    data['application/news-checkgroups'] = MimeType{'iana',[]string,false,''}
    data['application/news-groupinfo'] = MimeType{'iana',[]string,false,''}
    data['application/news-transmission'] = MimeType{'iana',[]string,false,''}
    data['application/nlsml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/node'] = MimeType{'iana',[]string,false,''}
    data['application/nss'] = MimeType{'iana',[]string,false,''}
    data['application/ocsp-request'] = MimeType{'iana',[]string,false,''}
    data['application/ocsp-response'] = MimeType{'iana',[]string,false,''}
    data['application/octet-stream'] = MimeType{'iana',['bin', 'dms', 'lrf', 'mar', 'so', 'dist', 'distz', 'pkg', 'bpk', 'dump', 'elc', 'deploy', 'exe', 'dll', 'deb', 'dmg', 'iso', 'img', 'msi', 'msp', 'msm', 'buffer'],false,''}
    data['application/oda'] = MimeType{'iana',['oda'],false,''}
    data['application/odm+xml'] = MimeType{'iana',[]string,true,''}
    data['application/odx'] = MimeType{'iana',[]string,false,''}
    data['application/oebps-package+xml'] = MimeType{'iana',['opf'],true,''}
    data['application/ogg'] = MimeType{'iana',['ogx'],false,''}
    data['application/omdoc+xml'] = MimeType{'apache',['omdoc'],true,''}
    data['application/onenote'] = MimeType{'apache',['onetoc', 'onetoc2', 'onetmp', 'onepkg'],false,''}
    data['application/oscore'] = MimeType{'iana',[]string,false,''}
    data['application/oxps'] = MimeType{'iana',['oxps'],false,''}
    data['application/p2p-overlay+xml'] = MimeType{'iana',[]string,true,''}
    data['application/parityfec'] = MimeType{'iana',[]string,false,''}
    data['application/passport'] = MimeType{'iana',[]string,false,''}
    data['application/patch-ops-error+xml'] = MimeType{'iana',['xer'],true,''}
    data['application/pdf'] = MimeType{'iana',['pdf'],false,''}
    data['application/pdx'] = MimeType{'iana',[]string,false,''}
    data['application/pem-certificate-chain'] = MimeType{'iana',[]string,false,''}
    data['application/pgp-encrypted'] = MimeType{'iana',['pgp'],false,''}
    data['application/pgp-keys'] = MimeType{'iana',[]string,false,''}
    data['application/pgp-signature'] = MimeType{'iana',['asc', 'sig'],false,''}
    data['application/pics-rules'] = MimeType{'apache',['prf'],false,''}
    data['application/pidf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/pidf-diff+xml'] = MimeType{'iana',[]string,true,''}
    data['application/pkcs10'] = MimeType{'iana',['p10'],false,''}
    data['application/pkcs12'] = MimeType{'iana',[]string,false,''}
    data['application/pkcs7-mime'] = MimeType{'iana',['p7m', 'p7c'],false,''}
    data['application/pkcs7-signature'] = MimeType{'iana',['p7s'],false,''}
    data['application/pkcs8'] = MimeType{'iana',['p8'],false,''}
    data['application/pkcs8-encrypted'] = MimeType{'iana',[]string,false,''}
    data['application/pkix-attr-cert'] = MimeType{'iana',['ac'],false,''}
    data['application/pkix-cert'] = MimeType{'iana',['cer'],false,''}
    data['application/pkix-crl'] = MimeType{'iana',['crl'],false,''}
    data['application/pkix-pkipath'] = MimeType{'iana',['pkipath'],false,''}
    data['application/pkixcmp'] = MimeType{'iana',['pki'],false,''}
    data['application/pls+xml'] = MimeType{'iana',['pls'],true,''}
    data['application/poc-settings+xml'] = MimeType{'iana',[]string,true,''}
    data['application/postscript'] = MimeType{'iana',['ai', 'eps', 'ps'],true,''}
    data['application/ppsp-tracker+json'] = MimeType{'iana',[]string,true,''}
    data['application/problem+json'] = MimeType{'iana',[]string,true,''}
    data['application/problem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/provenance+xml'] = MimeType{'iana',[]string,true,''}
    data['application/prs.alvestrand.titrax-sheet'] = MimeType{'iana',[]string,false,''}
    data['application/prs.cww'] = MimeType{'iana',['cww'],false,''}
    data['application/prs.hpub+zip'] = MimeType{'iana',[]string,false,''}
    data['application/prs.nprend'] = MimeType{'iana',[]string,false,''}
    data['application/prs.plucker'] = MimeType{'iana',[]string,false,''}
    data['application/prs.rdf-xml-crypt'] = MimeType{'iana',[]string,false,''}
    data['application/prs.xsf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/pskc+xml'] = MimeType{'iana',['pskcxml'],true,''}
    data['application/qsig'] = MimeType{'iana',[]string,false,''}
    data['application/raml+yaml'] = MimeType{'',['raml'],true,''}
    data['application/raptorfec'] = MimeType{'iana',[]string,false,''}
    data['application/rdap+json'] = MimeType{'iana',[]string,true,''}
    data['application/rdf+xml'] = MimeType{'iana',['rdf', 'owl'],true,''}
    data['application/reginfo+xml'] = MimeType{'iana',['rif'],true,''}
    data['application/relax-ng-compact-syntax'] = MimeType{'iana',['rnc'],false,''}
    data['application/remote-printing'] = MimeType{'iana',[]string,false,''}
    data['application/reputon+json'] = MimeType{'iana',[]string,true,''}
    data['application/resource-lists+xml'] = MimeType{'iana',['rl'],true,''}
    data['application/resource-lists-diff+xml'] = MimeType{'iana',['rld'],true,''}
    data['application/rfc+xml'] = MimeType{'iana',[]string,true,''}
    data['application/riscos'] = MimeType{'iana',[]string,false,''}
    data['application/rlmi+xml'] = MimeType{'iana',[]string,true,''}
    data['application/rls-services+xml'] = MimeType{'iana',['rs'],true,''}
    data['application/route-apd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/route-s-tsid+xml'] = MimeType{'iana',[]string,true,''}
    data['application/route-usd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/rpki-ghostbusters'] = MimeType{'iana',['gbr'],false,''}
    data['application/rpki-manifest'] = MimeType{'iana',['mft'],false,''}
    data['application/rpki-publication'] = MimeType{'iana',[]string,false,''}
    data['application/rpki-roa'] = MimeType{'iana',['roa'],false,''}
    data['application/rpki-updown'] = MimeType{'iana',[]string,false,''}
    data['application/rsd+xml'] = MimeType{'apache',['rsd'],true,''}
    data['application/rss+xml'] = MimeType{'apache',['rss'],true,''}
    data['application/rtf'] = MimeType{'iana',['rtf'],true,''}
    data['application/rtploopback'] = MimeType{'iana',[]string,false,''}
    data['application/rtx'] = MimeType{'iana',[]string,false,''}
    data['application/samlassertion+xml'] = MimeType{'iana',[]string,true,''}
    data['application/samlmetadata+xml'] = MimeType{'iana',[]string,true,''}
    data['application/sbml+xml'] = MimeType{'iana',['sbml'],true,''}
    data['application/scaip+xml'] = MimeType{'iana',[]string,true,''}
    data['application/scim+json'] = MimeType{'iana',[]string,true,''}
    data['application/scvp-cv-request'] = MimeType{'iana',['scq'],false,''}
    data['application/scvp-cv-response'] = MimeType{'iana',['scs'],false,''}
    data['application/scvp-vp-request'] = MimeType{'iana',['spq'],false,''}
    data['application/scvp-vp-response'] = MimeType{'iana',['spp'],false,''}
    data['application/sdp'] = MimeType{'iana',['sdp'],false,''}
    data['application/secevent+jwt'] = MimeType{'iana',[]string,false,''}
    data['application/senml+cbor'] = MimeType{'iana',[]string,false,''}
    data['application/senml+json'] = MimeType{'iana',[]string,true,''}
    data['application/senml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/senml-exi'] = MimeType{'iana',[]string,false,''}
    data['application/sensml+cbor'] = MimeType{'iana',[]string,false,''}
    data['application/sensml+json'] = MimeType{'iana',[]string,true,''}
    data['application/sensml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/sensml-exi'] = MimeType{'iana',[]string,false,''}
    data['application/sep+xml'] = MimeType{'iana',[]string,true,''}
    data['application/sep-exi'] = MimeType{'iana',[]string,false,''}
    data['application/session-info'] = MimeType{'iana',[]string,false,''}
    data['application/set-payment'] = MimeType{'iana',[]string,false,''}
    data['application/set-payment-initiation'] = MimeType{'iana',['setpay'],false,''}
    data['application/set-registration'] = MimeType{'iana',[]string,false,''}
    data['application/set-registration-initiation'] = MimeType{'iana',['setreg'],false,''}
    data['application/sgml'] = MimeType{'iana',[]string,false,''}
    data['application/sgml-open-catalog'] = MimeType{'iana',[]string,false,''}
    data['application/shf+xml'] = MimeType{'iana',['shf'],true,''}
    data['application/sieve'] = MimeType{'iana',['siv', 'sieve'],false,''}
    data['application/simple-filter+xml'] = MimeType{'iana',[]string,true,''}
    data['application/simple-message-summary'] = MimeType{'iana',[]string,false,''}
    data['application/simplesymbolcontainer'] = MimeType{'iana',[]string,false,''}
    data['application/slate'] = MimeType{'iana',[]string,false,''}
    data['application/smil'] = MimeType{'iana',[]string,false,''}
    data['application/smil+xml'] = MimeType{'iana',['smi', 'smil'],true,''}
    data['application/smpte336m'] = MimeType{'iana',[]string,false,''}
    data['application/soap+fastinfoset'] = MimeType{'iana',[]string,false,''}
    data['application/soap+xml'] = MimeType{'iana',[]string,true,''}
    data['application/sparql-query'] = MimeType{'iana',['rq'],false,''}
    data['application/sparql-results+xml'] = MimeType{'iana',['srx'],true,''}
    data['application/spirits-event+xml'] = MimeType{'iana',[]string,true,''}
    data['application/sql'] = MimeType{'iana',[]string,false,''}
    data['application/srgs'] = MimeType{'iana',['gram'],false,''}
    data['application/srgs+xml'] = MimeType{'iana',['grxml'],true,''}
    data['application/sru+xml'] = MimeType{'iana',['sru'],true,''}
    data['application/ssdl+xml'] = MimeType{'apache',['ssdl'],true,''}
    data['application/ssml+xml'] = MimeType{'iana',['ssml'],true,''}
    data['application/stix+json'] = MimeType{'iana',[]string,true,''}
    data['application/tamp-apex-update'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-apex-update-confirm'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-community-update'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-community-update-confirm'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-error'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-sequence-adjust'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-sequence-adjust-confirm'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-status-query'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-status-response'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-update'] = MimeType{'iana',[]string,false,''}
    data['application/tamp-update-confirm'] = MimeType{'iana',[]string,false,''}
    data['application/tar'] = MimeType{'',[]string,true,''}
    data['application/taxii+json'] = MimeType{'iana',[]string,true,''}
    data['application/tei+xml'] = MimeType{'iana',['tei', 'teicorpus'],true,''}
    data['application/tetra_isi'] = MimeType{'iana',[]string,false,''}
    data['application/thraud+xml'] = MimeType{'iana',['tfi'],true,''}
    data['application/timestamp-query'] = MimeType{'iana',[]string,false,''}
    data['application/timestamp-reply'] = MimeType{'iana',[]string,false,''}
    data['application/timestamped-data'] = MimeType{'iana',['tsd'],false,''}
    data['application/tlsrpt+gzip'] = MimeType{'iana',[]string,false,''}
    data['application/tlsrpt+json'] = MimeType{'iana',[]string,true,''}
    data['application/tnauthlist'] = MimeType{'iana',[]string,false,''}
    data['application/trickle-ice-sdpfrag'] = MimeType{'iana',[]string,false,''}
    data['application/trig'] = MimeType{'iana',[]string,false,''}
    data['application/ttml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/tve-trigger'] = MimeType{'iana',[]string,false,''}
    data['application/tzif'] = MimeType{'iana',[]string,false,''}
    data['application/tzif-leap'] = MimeType{'iana',[]string,false,''}
    data['application/ulpfec'] = MimeType{'iana',[]string,false,''}
    data['application/urc-grpsheet+xml'] = MimeType{'iana',[]string,true,''}
    data['application/urc-ressheet+xml'] = MimeType{'iana',[]string,true,''}
    data['application/urc-targetdesc+xml'] = MimeType{'iana',[]string,true,''}
    data['application/urc-uisocketdesc+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vcard+json'] = MimeType{'iana',[]string,true,''}
    data['application/vcard+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vemmi'] = MimeType{'iana',[]string,false,''}
    data['application/vividence.scriptfile'] = MimeType{'apache',[]string,false,''}
    data['application/vnd.1000minds.decision-model+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp-prose+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp-prose-pc3ch+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp-v2x-local-service-information'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3gpp.access-transfer-events+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.bsf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.gmop+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mc-signalling-ear'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3gpp.mcdata-affiliation-command+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcdata-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcdata-payload'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3gpp.mcdata-service-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcdata-signalling'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3gpp.mcdata-ue-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcdata-user-profile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-affiliation-command+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-floor-request+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-location-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-mbms-usage-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-service-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-signed+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-ue-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-ue-init-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcptt-user-profile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-affiliation-command+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-affiliation-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-location-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-mbms-usage-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-service-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-transmission-request+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-ue-config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mcvideo-user-profile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.mid-call+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.pic-bw-large'] = MimeType{'iana',['plb'],false,''}
    data['application/vnd.3gpp.pic-bw-small'] = MimeType{'iana',['psb'],false,''}
    data['application/vnd.3gpp.pic-bw-var'] = MimeType{'iana',['pvb'],false,''}
    data['application/vnd.3gpp.sms'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3gpp.sms+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.srvcc-ext+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.srvcc-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.state-and-event-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp.ussd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp2.bcmcsinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.3gpp2.sms'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3gpp2.tcap'] = MimeType{'iana',['tcap'],false,''}
    data['application/vnd.3lightssoftware.imagescal'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.3m.post-it-notes'] = MimeType{'iana',['pwn'],false,''}
    data['application/vnd.accpac.simply.aso'] = MimeType{'iana',['aso'],false,''}
    data['application/vnd.accpac.simply.imp'] = MimeType{'iana',['imp'],false,''}
    data['application/vnd.acucobol'] = MimeType{'iana',['acu'],false,''}
    data['application/vnd.acucorp'] = MimeType{'iana',['atc', 'acutc'],false,''}
    data['application/vnd.adobe.air-application-installer-package+zip'] = MimeType{'apache',['air'],false,''}
    data['application/vnd.adobe.flash.movie'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.adobe.formscentral.fcdt'] = MimeType{'iana',['fcdt'],false,''}
    data['application/vnd.adobe.fxp'] = MimeType{'iana',['fxp', 'fxpl'],false,''}
    data['application/vnd.adobe.partial-upload'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.adobe.xdp+xml'] = MimeType{'iana',['xdp'],true,''}
    data['application/vnd.adobe.xfdf'] = MimeType{'iana',['xfdf'],false,''}
    data['application/vnd.aether.imp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.afpc.afplinedata'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.afpc.modca'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ah-barcode'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ahead.space'] = MimeType{'iana',['ahead'],false,''}
    data['application/vnd.airzip.filesecure.azf'] = MimeType{'iana',['azf'],false,''}
    data['application/vnd.airzip.filesecure.azs'] = MimeType{'iana',['azs'],false,''}
    data['application/vnd.amadeus+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.amazon.ebook'] = MimeType{'apache',['azw'],false,''}
    data['application/vnd.amazon.mobi8-ebook'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.americandynamics.acc'] = MimeType{'iana',['acc'],false,''}
    data['application/vnd.amiga.ami'] = MimeType{'iana',['ami'],false,''}
    data['application/vnd.amundsen.maze+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.android.package-archive'] = MimeType{'apache',['apk'],false,''}
    data['application/vnd.anki'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.anser-web-certificate-issue-initiation'] = MimeType{'iana',['cii'],false,''}
    data['application/vnd.anser-web-funds-transfer-initiation'] = MimeType{'apache',['fti'],false,''}
    data['application/vnd.antix.game-component'] = MimeType{'iana',['atx'],false,''}
    data['application/vnd.apache.thrift.binary'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.apache.thrift.compact'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.apache.thrift.json'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.api+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.apothekende.reservation+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.apple.installer+xml'] = MimeType{'iana',['mpkg'],true,''}
    data['application/vnd.apple.keynote'] = MimeType{'iana',['keynote'],false,''}
    data['application/vnd.apple.mpegurl'] = MimeType{'iana',['m3u8'],false,''}
    data['application/vnd.apple.numbers'] = MimeType{'iana',['numbers'],false,''}
    data['application/vnd.apple.pages'] = MimeType{'iana',['pages'],false,''}
    data['application/vnd.apple.pkpass'] = MimeType{'',['pkpass'],false,''}
    data['application/vnd.arastra.swi'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.aristanetworks.swi'] = MimeType{'iana',['swi'],false,''}
    data['application/vnd.artisan+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.artsquare'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.astraea-software.iota'] = MimeType{'iana',['iota'],false,''}
    data['application/vnd.audiograph'] = MimeType{'iana',['aep'],false,''}
    data['application/vnd.autopackage'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.avalon+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.avistar+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.balsamiq.bmml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.balsamiq.bmpr'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.banana-accounting'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.bbf.usp.msg'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.bbf.usp.msg+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.bekitzur-stech+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.bint.med-content'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.biopax.rdf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.blink-idb-value-wrapper'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.blueice.multipass'] = MimeType{'iana',['mpm'],false,''}
    data['application/vnd.bluetooth.ep.oob'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.bluetooth.le.oob'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.bmi'] = MimeType{'iana',['bmi'],false,''}
    data['application/vnd.businessobjects'] = MimeType{'iana',['rep'],false,''}
    data['application/vnd.byu.uapi+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.cab-jscript'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.canon-cpdl'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.canon-lips'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.capasystems-pg+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.cendio.thinlinc.clientconf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.century-systems.tcp_stream'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.chemdraw+xml'] = MimeType{'iana',['cdxml'],true,''}
    data['application/vnd.chess-pgn'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.chipnuts.karaoke-mmd'] = MimeType{'iana',['mmd'],false,''}
    data['application/vnd.cinderella'] = MimeType{'iana',['cdy'],false,''}
    data['application/vnd.cirpack.isdn-ext'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.citationstyles.style+xml'] = MimeType{'iana',['csl'],true,''}
    data['application/vnd.claymore'] = MimeType{'iana',['cla'],false,''}
    data['application/vnd.cloanto.rp9'] = MimeType{'iana',['rp9'],false,''}
    data['application/vnd.clonk.c4group'] = MimeType{'iana',['c4g', 'c4d', 'c4f', 'c4p', 'c4u'],false,''}
    data['application/vnd.cluetrust.cartomobile-config'] = MimeType{'iana',['c11amc'],false,''}
    data['application/vnd.cluetrust.cartomobile-config-pkg'] = MimeType{'iana',['c11amz'],false,''}
    data['application/vnd.coffeescript'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collabio.xodocuments.document'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collabio.xodocuments.document-template'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collabio.xodocuments.presentation'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collabio.xodocuments.presentation-template'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collabio.xodocuments.spreadsheet'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collabio.xodocuments.spreadsheet-template'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.collection+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.collection.doc+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.collection.next+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.comicbook+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.comicbook-rar'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.commerce-battelle'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.commonspace'] = MimeType{'iana',['csp'],false,''}
    data['application/vnd.contact.cmsg'] = MimeType{'iana',['cdbcmsg'],false,''}
    data['application/vnd.coreos.ignition+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.cosmocaller'] = MimeType{'iana',['cmc'],false,''}
    data['application/vnd.crick.clicker'] = MimeType{'iana',['clkx'],false,''}
    data['application/vnd.crick.clicker.keyboard'] = MimeType{'iana',['clkk'],false,''}
    data['application/vnd.crick.clicker.palette'] = MimeType{'iana',['clkp'],false,''}
    data['application/vnd.crick.clicker.template'] = MimeType{'iana',['clkt'],false,''}
    data['application/vnd.crick.clicker.wordbank'] = MimeType{'iana',['clkw'],false,''}
    data['application/vnd.criticaltools.wbs+xml'] = MimeType{'iana',['wbs'],true,''}
    data['application/vnd.ctc-posml'] = MimeType{'iana',['pml'],false,''}
    data['application/vnd.ctct.ws+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.cups-pdf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.cups-postscript'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.cups-ppd'] = MimeType{'iana',['ppd'],false,''}
    data['application/vnd.cups-raster'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.cups-raw'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.curl'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.curl.car'] = MimeType{'apache',['car'],false,''}
    data['application/vnd.curl.pcurl'] = MimeType{'apache',['pcurl'],false,''}
    data['application/vnd.cyan.dean.root+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.cybank'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.d2l.coursepackage1p0+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dart'] = MimeType{'iana',['dart'],true,''}
    data['application/vnd.data-vision.rdz'] = MimeType{'iana',['rdz'],false,''}
    data['application/vnd.datapackage+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dataresource+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.debian.binary-package'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dece.data'] = MimeType{'iana',['uvf', 'uvvf', 'uvd', 'uvvd'],false,''}
    data['application/vnd.dece.ttml+xml'] = MimeType{'iana',['uvt', 'uvvt'],true,''}
    data['application/vnd.dece.unspecified'] = MimeType{'iana',['uvx', 'uvvx'],false,''}
    data['application/vnd.dece.zip'] = MimeType{'iana',['uvz', 'uvvz'],false,''}
    data['application/vnd.denovo.fcselayout-link'] = MimeType{'iana',['fe_launch'],false,''}
    data['application/vnd.desmume.movie'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dir-bi.plate-dl-nosuffix'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dm.delegation+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dna'] = MimeType{'iana',['dna'],false,''}
    data['application/vnd.document+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dolby.mlp'] = MimeType{'apache',['mlp'],false,''}
    data['application/vnd.dolby.mobile.1'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dolby.mobile.2'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.doremir.scorecloud-binary-document'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dpgraph'] = MimeType{'iana',['dpg'],false,''}
    data['application/vnd.dreamfactory'] = MimeType{'iana',['dfac'],false,''}
    data['application/vnd.drive+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ds-keypoint'] = MimeType{'apache',['kpxx'],false,''}
    data['application/vnd.dtg.local'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dtg.local.flash'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dtg.local.html'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.ait'] = MimeType{'iana',['ait'],false,''}
    data['application/vnd.dvb.dvbj'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.esgcontainer'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.ipdcdftnotifaccess'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.ipdcesgaccess'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.ipdcesgaccess2'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.ipdcesgpdd'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.ipdcroaming'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.iptv.alfec-base'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.iptv.alfec-enhancement'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.notif-aggregate-root+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.notif-container+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.notif-generic+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.notif-ia-msglist+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.notif-ia-registration-request+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.notif-ia-registration-response+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.notif-init+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.dvb.pfr'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dvb.service'] = MimeType{'iana',['svc'],false,''}
    data['application/vnd.dxr'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.dynageo'] = MimeType{'iana',['geo'],false,''}
    data['application/vnd.dzr'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.easykaraoke.cdgdownload'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecdis-update'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecip.rlp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecowin.chart'] = MimeType{'iana',['mag'],false,''}
    data['application/vnd.ecowin.filerequest'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecowin.fileupdate'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecowin.series'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecowin.seriesrequest'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ecowin.seriesupdate'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.efi.img'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.efi.iso'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.emclient.accessrequest+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.enliven'] = MimeType{'iana',['nml'],false,''}
    data['application/vnd.enphase.envoy'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.eprints.data+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.epson.esf'] = MimeType{'iana',['esf'],false,''}
    data['application/vnd.epson.msf'] = MimeType{'iana',['msf'],false,''}
    data['application/vnd.epson.quickanime'] = MimeType{'iana',['qam'],false,''}
    data['application/vnd.epson.salt'] = MimeType{'iana',['slt'],false,''}
    data['application/vnd.epson.ssf'] = MimeType{'iana',['ssf'],false,''}
    data['application/vnd.ericsson.quickcall'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.espass-espass+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.eszigno3+xml'] = MimeType{'iana',['es3', 'et3'],true,''}
    data['application/vnd.etsi.aoc+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.asic-e+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.etsi.asic-s+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.etsi.cug+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvcommand+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvdiscovery+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvprofile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvsad-bc+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvsad-cod+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvsad-npvr+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvservice+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvsync+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.iptvueprofile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.mcid+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.mheg5'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.etsi.overload-control-policy-dataset+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.pstn+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.sci+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.simservs+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.timestamp-token'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.etsi.tsl+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.etsi.tsl.der'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.eudora.data'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.evolv.ecig.profile'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.evolv.ecig.settings'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.evolv.ecig.theme'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.exstream-empower+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.exstream-package'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ezpix-album'] = MimeType{'iana',['ez2'],false,''}
    data['application/vnd.ezpix-package'] = MimeType{'iana',['ez3'],false,''}
    data['application/vnd.f-secure.mobile'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fastcopy-disk-image'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fdf'] = MimeType{'iana',['fdf'],false,''}
    data['application/vnd.fdsn.mseed'] = MimeType{'iana',['mseed'],false,''}
    data['application/vnd.fdsn.seed'] = MimeType{'iana',['seed', 'dataless'],false,''}
    data['application/vnd.ffsns'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.filmit.zfc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fints'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.firemonkeys.cloudcell'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.flographit'] = MimeType{'iana',['gph'],false,''}
    data['application/vnd.fluxtime.clip'] = MimeType{'iana',['ftc'],false,''}
    data['application/vnd.font-fontforge-sfd'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.framemaker'] = MimeType{'iana',['fm', 'frame', 'maker', 'book'],false,''}
    data['application/vnd.frogans.fnc'] = MimeType{'iana',['fnc'],false,''}
    data['application/vnd.frogans.ltf'] = MimeType{'iana',['ltf'],false,''}
    data['application/vnd.fsc.weblaunch'] = MimeType{'iana',['fsc'],false,''}
    data['application/vnd.fujitsu.oasys'] = MimeType{'iana',['oas'],false,''}
    data['application/vnd.fujitsu.oasys2'] = MimeType{'iana',['oa2'],false,''}
    data['application/vnd.fujitsu.oasys3'] = MimeType{'iana',['oa3'],false,''}
    data['application/vnd.fujitsu.oasysgp'] = MimeType{'iana',['fg5'],false,''}
    data['application/vnd.fujitsu.oasysprs'] = MimeType{'iana',['bh2'],false,''}
    data['application/vnd.fujixerox.art-ex'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fujixerox.art4'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fujixerox.ddd'] = MimeType{'iana',['ddd'],false,''}
    data['application/vnd.fujixerox.docuworks'] = MimeType{'iana',['xdw'],false,''}
    data['application/vnd.fujixerox.docuworks.binder'] = MimeType{'iana',['xbd'],false,''}
    data['application/vnd.fujixerox.docuworks.container'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fujixerox.hbpl'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.fut-misnet'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.futoin+cbor'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.futoin+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.fuzzysheet'] = MimeType{'iana',['fzs'],false,''}
    data['application/vnd.genomatix.tuxedo'] = MimeType{'iana',['txd'],false,''}
    data['application/vnd.geo+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.geocube+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.geogebra.file'] = MimeType{'iana',['ggb'],false,''}
    data['application/vnd.geogebra.tool'] = MimeType{'iana',['ggt'],false,''}
    data['application/vnd.geometry-explorer'] = MimeType{'iana',['gex', 'gre'],false,''}
    data['application/vnd.geonext'] = MimeType{'iana',['gxt'],false,''}
    data['application/vnd.geoplan'] = MimeType{'iana',['g2w'],false,''}
    data['application/vnd.geospace'] = MimeType{'iana',['g3w'],false,''}
    data['application/vnd.gerber'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.globalplatform.card-content-mgt'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.globalplatform.card-content-mgt-response'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.gmx'] = MimeType{'iana',['gmx'],false,''}
    data['application/vnd.google-apps.document'] = MimeType{'',['gdoc'],false,''}
    data['application/vnd.google-apps.presentation'] = MimeType{'',['gslides'],false,''}
    data['application/vnd.google-apps.spreadsheet'] = MimeType{'',['gsheet'],false,''}
    data['application/vnd.google-earth.kml+xml'] = MimeType{'iana',['kml'],true,''}
    data['application/vnd.google-earth.kmz'] = MimeType{'iana',['kmz'],false,''}
    data['application/vnd.gov.sk.e-form+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.gov.sk.e-form+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.gov.sk.xmldatacontainer+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.grafeq'] = MimeType{'iana',['gqf', 'gqs'],false,''}
    data['application/vnd.gridmp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.groove-account'] = MimeType{'iana',['gac'],false,''}
    data['application/vnd.groove-help'] = MimeType{'iana',['ghf'],false,''}
    data['application/vnd.groove-identity-message'] = MimeType{'iana',['gim'],false,''}
    data['application/vnd.groove-injector'] = MimeType{'iana',['grv'],false,''}
    data['application/vnd.groove-tool-message'] = MimeType{'iana',['gtm'],false,''}
    data['application/vnd.groove-tool-template'] = MimeType{'iana',['tpl'],false,''}
    data['application/vnd.groove-vcard'] = MimeType{'iana',['vcg'],false,''}
    data['application/vnd.hal+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.hal+xml'] = MimeType{'iana',['hal'],true,''}
    data['application/vnd.handheld-entertainment+xml'] = MimeType{'iana',['zmm'],true,''}
    data['application/vnd.hbci'] = MimeType{'iana',['hbci'],false,''}
    data['application/vnd.hc+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.hcl-bireports'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.hdt'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.heroku+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.hhe.lesson-player'] = MimeType{'iana',['les'],false,''}
    data['application/vnd.hp-hpgl'] = MimeType{'iana',['hpgl'],false,''}
    data['application/vnd.hp-hpid'] = MimeType{'iana',['hpid'],false,''}
    data['application/vnd.hp-hps'] = MimeType{'iana',['hps'],false,''}
    data['application/vnd.hp-jlyt'] = MimeType{'iana',['jlt'],false,''}
    data['application/vnd.hp-pcl'] = MimeType{'iana',['pcl'],false,''}
    data['application/vnd.hp-pclxl'] = MimeType{'iana',['pclxl'],false,''}
    data['application/vnd.httphone'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.hydrostatix.sof-data'] = MimeType{'iana',['sfd-hdstx'],false,''}
    data['application/vnd.hyper+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.hyper-item+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.hyperdrive+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.hzn-3d-crossword'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ibm.afplinedata'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ibm.electronic-media'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ibm.minipay'] = MimeType{'iana',['mpy'],false,''}
    data['application/vnd.ibm.modcap'] = MimeType{'iana',['afp', 'listafp', 'list3820'],false,''}
    data['application/vnd.ibm.rights-management'] = MimeType{'iana',['irm'],false,''}
    data['application/vnd.ibm.secure-container'] = MimeType{'iana',['sc'],false,''}
    data['application/vnd.iccprofile'] = MimeType{'iana',['icc', 'icm'],false,''}
    data['application/vnd.ieee.1905'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.igloader'] = MimeType{'iana',['igl'],false,''}
    data['application/vnd.imagemeter.folder+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.imagemeter.image+zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.immervision-ivp'] = MimeType{'iana',['ivp'],false,''}
    data['application/vnd.immervision-ivu'] = MimeType{'iana',['ivu'],false,''}
    data['application/vnd.ims.imsccv1p1'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ims.imsccv1p2'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ims.imsccv1p3'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ims.lis.v2.result+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ims.lti.v2.toolconsumerprofile+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ims.lti.v2.toolproxy+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ims.lti.v2.toolproxy.id+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ims.lti.v2.toolsettings+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ims.lti.v2.toolsettings.simple+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.informedcontrol.rms+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.informix-visionary'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.infotech.project'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.infotech.project+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.innopath.wamp.notification'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.insors.igm'] = MimeType{'iana',['igm'],false,''}
    data['application/vnd.intercon.formnet'] = MimeType{'iana',['xpw', 'xpx'],false,''}
    data['application/vnd.intergeo'] = MimeType{'iana',['i2g'],false,''}
    data['application/vnd.intertrust.digibox'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.intertrust.nncp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.intu.qbo'] = MimeType{'iana',['qbo'],false,''}
    data['application/vnd.intu.qfx'] = MimeType{'iana',['qfx'],false,''}
    data['application/vnd.iptc.g2.catalogitem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.iptc.g2.conceptitem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.iptc.g2.knowledgeitem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.iptc.g2.newsitem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.iptc.g2.newsmessage+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.iptc.g2.packageitem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.iptc.g2.planningitem+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ipunplugged.rcprofile'] = MimeType{'iana',['rcprofile'],false,''}
    data['application/vnd.irepository.package+xml'] = MimeType{'iana',['irp'],true,''}
    data['application/vnd.is-xpr'] = MimeType{'iana',['xpr'],false,''}
    data['application/vnd.isac.fcs'] = MimeType{'iana',['fcs'],false,''}
    data['application/vnd.jam'] = MimeType{'iana',['jam'],false,''}
    data['application/vnd.japannet-directory-service'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-jpnstore-wakeup'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-payment-wakeup'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-registration'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-registration-wakeup'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-setstore-wakeup'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-verification'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.japannet-verification-wakeup'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.jcp.javame.midlet-rms'] = MimeType{'iana',['rms'],false,''}
    data['application/vnd.jisp'] = MimeType{'iana',['jisp'],false,''}
    data['application/vnd.joost.joda-archive'] = MimeType{'iana',['joda'],false,''}
    data['application/vnd.jsk.isdn-ngn'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.kahootz'] = MimeType{'iana',['ktz', 'ktr'],false,''}
    data['application/vnd.kde.karbon'] = MimeType{'iana',['karbon'],false,''}
    data['application/vnd.kde.kchart'] = MimeType{'iana',['chrt'],false,''}
    data['application/vnd.kde.kformula'] = MimeType{'iana',['kfo'],false,''}
    data['application/vnd.kde.kivio'] = MimeType{'iana',['flw'],false,''}
    data['application/vnd.kde.kontour'] = MimeType{'iana',['kon'],false,''}
    data['application/vnd.kde.kpresenter'] = MimeType{'iana',['kpr', 'kpt'],false,''}
    data['application/vnd.kde.kspread'] = MimeType{'iana',['ksp'],false,''}
    data['application/vnd.kde.kword'] = MimeType{'iana',['kwd', 'kwt'],false,''}
    data['application/vnd.kenameaapp'] = MimeType{'iana',['htke'],false,''}
    data['application/vnd.kidspiration'] = MimeType{'iana',['kia'],false,''}
    data['application/vnd.kinar'] = MimeType{'iana',['kne', 'knp'],false,''}
    data['application/vnd.koan'] = MimeType{'iana',['skp', 'skd', 'skt', 'skm'],false,''}
    data['application/vnd.kodak-descriptor'] = MimeType{'iana',['sse'],false,''}
    data['application/vnd.las.las+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.las.las+xml'] = MimeType{'iana',['lasxml'],true,''}
    data['application/vnd.leap+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.liberty-request+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.llamagraphics.life-balance.desktop'] = MimeType{'iana',['lbd'],false,''}
    data['application/vnd.llamagraphics.life-balance.exchange+xml'] = MimeType{'iana',['lbe'],true,''}
    data['application/vnd.lotus-1-2-3'] = MimeType{'iana',['123'],false,''}
    data['application/vnd.lotus-approach'] = MimeType{'iana',['apr'],false,''}
    data['application/vnd.lotus-freelance'] = MimeType{'iana',['pre'],false,''}
    data['application/vnd.lotus-notes'] = MimeType{'iana',['nsf'],false,''}
    data['application/vnd.lotus-organizer'] = MimeType{'iana',['org'],false,''}
    data['application/vnd.lotus-screencam'] = MimeType{'iana',['scm'],false,''}
    data['application/vnd.lotus-wordpro'] = MimeType{'iana',['lwp'],false,''}
    data['application/vnd.macports.portpkg'] = MimeType{'iana',['portpkg'],false,''}
    data['application/vnd.mapbox-vector-tile'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.marlin.drm.actiontoken+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.marlin.drm.conftoken+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.marlin.drm.license+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.marlin.drm.mdcf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mason+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.maxmind.maxmind-db'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mcd'] = MimeType{'iana',['mcd'],false,''}
    data['application/vnd.medcalcdata'] = MimeType{'iana',['mc1'],false,''}
    data['application/vnd.mediastation.cdkey'] = MimeType{'iana',['cdkey'],false,''}
    data['application/vnd.meridian-slingshot'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mfer'] = MimeType{'iana',['mwf'],false,''}
    data['application/vnd.mfmp'] = MimeType{'iana',['mfm'],false,''}
    data['application/vnd.micro+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.micrografx.flo'] = MimeType{'iana',['flo'],false,''}
    data['application/vnd.micrografx.igx'] = MimeType{'iana',['igx'],false,''}
    data['application/vnd.microsoft.portable-executable'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.microsoft.windows.thumbnail-cache'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.miele+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.mif'] = MimeType{'iana',['mif'],false,''}
    data['application/vnd.minisoft-hp3000-save'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mitsubishi.misty-guard.trustweb'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mobius.daf'] = MimeType{'iana',['daf'],false,''}
    data['application/vnd.mobius.dis'] = MimeType{'iana',['dis'],false,''}
    data['application/vnd.mobius.mbk'] = MimeType{'iana',['mbk'],false,''}
    data['application/vnd.mobius.mqy'] = MimeType{'iana',['mqy'],false,''}
    data['application/vnd.mobius.msl'] = MimeType{'iana',['msl'],false,''}
    data['application/vnd.mobius.plc'] = MimeType{'iana',['plc'],false,''}
    data['application/vnd.mobius.txf'] = MimeType{'iana',['txf'],false,''}
    data['application/vnd.mophun.application'] = MimeType{'iana',['mpn'],false,''}
    data['application/vnd.mophun.certificate'] = MimeType{'iana',['mpc'],false,''}
    data['application/vnd.motorola.flexsuite'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.flexsuite.adsi'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.flexsuite.fis'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.flexsuite.gotap'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.flexsuite.kmr'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.flexsuite.ttc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.flexsuite.wem'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.motorola.iprm'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mozilla.xul+xml'] = MimeType{'iana',['xul'],true,''}
    data['application/vnd.ms-3mfdocument'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-artgalry'] = MimeType{'iana',['cil'],false,''}
    data['application/vnd.ms-asf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-cab-compressed'] = MimeType{'iana',['cab'],false,''}
    data['application/vnd.ms-color.iccprofile'] = MimeType{'apache',[]string,false,''}
    data['application/vnd.ms-excel'] = MimeType{'iana',['xls', 'xlm', 'xla', 'xlc', 'xlt', 'xlw'],false,''}
    data['application/vnd.ms-excel.addin.macroenabled.12'] = MimeType{'iana',['xlam'],false,''}
    data['application/vnd.ms-excel.sheet.binary.macroenabled.12'] = MimeType{'iana',['xlsb'],false,''}
    data['application/vnd.ms-excel.sheet.macroenabled.12'] = MimeType{'iana',['xlsm'],false,''}
    data['application/vnd.ms-excel.template.macroenabled.12'] = MimeType{'iana',['xltm'],false,''}
    data['application/vnd.ms-fontobject'] = MimeType{'iana',['eot'],true,''}
    data['application/vnd.ms-htmlhelp'] = MimeType{'iana',['chm'],false,''}
    data['application/vnd.ms-ims'] = MimeType{'iana',['ims'],false,''}
    data['application/vnd.ms-lrm'] = MimeType{'iana',['lrm'],false,''}
    data['application/vnd.ms-office.activex+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ms-officetheme'] = MimeType{'iana',['thmx'],false,''}
    data['application/vnd.ms-opentype'] = MimeType{'apache',[]string,true,''}
    data['application/vnd.ms-outlook'] = MimeType{'',['msg'],false,''}
    data['application/vnd.ms-package.obfuscated-opentype'] = MimeType{'apache',[]string,false,''}
    data['application/vnd.ms-pki.seccat'] = MimeType{'apache',['cat'],false,''}
    data['application/vnd.ms-pki.stl'] = MimeType{'apache',['stl'],false,''}
    data['application/vnd.ms-playready.initiator+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ms-powerpoint'] = MimeType{'iana',['ppt', 'pps', 'pot'],false,''}
    data['application/vnd.ms-powerpoint.addin.macroenabled.12'] = MimeType{'iana',['ppam'],false,''}
    data['application/vnd.ms-powerpoint.presentation.macroenabled.12'] = MimeType{'iana',['pptm'],false,''}
    data['application/vnd.ms-powerpoint.slide.macroenabled.12'] = MimeType{'iana',['sldm'],false,''}
    data['application/vnd.ms-powerpoint.slideshow.macroenabled.12'] = MimeType{'iana',['ppsm'],false,''}
    data['application/vnd.ms-powerpoint.template.macroenabled.12'] = MimeType{'iana',['potm'],false,''}
    data['application/vnd.ms-printdevicecapabilities+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ms-printing.printticket+xml'] = MimeType{'apache',[]string,true,''}
    data['application/vnd.ms-printschematicket+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.ms-project'] = MimeType{'iana',['mpp', 'mpt'],false,''}
    data['application/vnd.ms-tnef'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-windows.devicepairing'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-windows.nwprinting.oob'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-windows.printerpairing'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-windows.wsd.oob'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-wmdrm.lic-chlg-req'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-wmdrm.lic-resp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-wmdrm.meter-chlg-req'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-wmdrm.meter-resp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ms-word.document.macroenabled.12'] = MimeType{'iana',['docm'],false,''}
    data['application/vnd.ms-word.template.macroenabled.12'] = MimeType{'iana',['dotm'],false,''}
    data['application/vnd.ms-works'] = MimeType{'iana',['wps', 'wks', 'wcm', 'wdb'],false,''}
    data['application/vnd.ms-wpl'] = MimeType{'iana',['wpl'],false,''}
    data['application/vnd.ms-xpsdocument'] = MimeType{'iana',['xps'],false,''}
    data['application/vnd.msa-disk-image'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.mseq'] = MimeType{'iana',['mseq'],false,''}
    data['application/vnd.msign'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.multiad.creator'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.multiad.creator.cif'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.music-niff'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.musician'] = MimeType{'iana',['mus'],false,''}
    data['application/vnd.muvee.style'] = MimeType{'iana',['msty'],false,''}
    data['application/vnd.mynfc'] = MimeType{'iana',['taglet'],false,''}
    data['application/vnd.ncd.control'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ncd.reference'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nearst.inv+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nervana'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.netfpx'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.neurolanguage.nlu'] = MimeType{'iana',['nlu'],false,''}
    data['application/vnd.nimn'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nintendo.nitro.rom'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nintendo.snes.rom'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nitf'] = MimeType{'iana',['ntf', 'nitf'],false,''}
    data['application/vnd.noblenet-directory'] = MimeType{'iana',['nnd'],false,''}
    data['application/vnd.noblenet-sealer'] = MimeType{'iana',['nns'],false,''}
    data['application/vnd.noblenet-web'] = MimeType{'iana',['nnw'],false,''}
    data['application/vnd.nokia.catalogs'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nokia.conml+wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nokia.conml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nokia.iptv.config+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nokia.isds-radio-presets'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nokia.landmark+wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nokia.landmark+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nokia.landmarkcollection+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nokia.n-gage.ac+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nokia.n-gage.data'] = MimeType{'iana',['ngdat'],false,''}
    data['application/vnd.nokia.n-gage.symbian.install'] = MimeType{'iana',['n-gage'],false,''}
    data['application/vnd.nokia.ncd'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nokia.pcd+wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.nokia.pcd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.nokia.radio-preset'] = MimeType{'iana',['rpst'],false,''}
    data['application/vnd.nokia.radio-presets'] = MimeType{'iana',['rpss'],false,''}
    data['application/vnd.novadigm.edm'] = MimeType{'iana',['edm'],false,''}
    data['application/vnd.novadigm.edx'] = MimeType{'iana',['edx'],false,''}
    data['application/vnd.novadigm.ext'] = MimeType{'iana',['ext'],false,''}
    data['application/vnd.ntt-local.content-share'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ntt-local.file-transfer'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ntt-local.ogw_remote-access'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ntt-local.sip-ta_remote'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ntt-local.sip-ta_tcp_stream'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oasis.opendocument.chart'] = MimeType{'iana',['odc'],false,''}
    data['application/vnd.oasis.opendocument.chart-template'] = MimeType{'iana',['otc'],false,''}
    data['application/vnd.oasis.opendocument.database'] = MimeType{'iana',['odb'],false,''}
    data['application/vnd.oasis.opendocument.formula'] = MimeType{'iana',['odf'],false,''}
    data['application/vnd.oasis.opendocument.formula-template'] = MimeType{'iana',['odft'],false,''}
    data['application/vnd.oasis.opendocument.graphics'] = MimeType{'iana',['odg'],false,''}
    data['application/vnd.oasis.opendocument.graphics-template'] = MimeType{'iana',['otg'],false,''}
    data['application/vnd.oasis.opendocument.image'] = MimeType{'iana',['odi'],false,''}
    data['application/vnd.oasis.opendocument.image-template'] = MimeType{'iana',['oti'],false,''}
    data['application/vnd.oasis.opendocument.presentation'] = MimeType{'iana',['odp'],false,''}
    data['application/vnd.oasis.opendocument.presentation-template'] = MimeType{'iana',['otp'],false,''}
    data['application/vnd.oasis.opendocument.spreadsheet'] = MimeType{'iana',['ods'],false,''}
    data['application/vnd.oasis.opendocument.spreadsheet-template'] = MimeType{'iana',['ots'],false,''}
    data['application/vnd.oasis.opendocument.text'] = MimeType{'iana',['odt'],false,''}
    data['application/vnd.oasis.opendocument.text-master'] = MimeType{'iana',['odm'],false,''}
    data['application/vnd.oasis.opendocument.text-template'] = MimeType{'iana',['ott'],false,''}
    data['application/vnd.oasis.opendocument.text-web'] = MimeType{'iana',['oth'],false,''}
    data['application/vnd.obn'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ocf+cbor'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oftn.l10n+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.contentaccessdownload+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.contentaccessstreaming+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.cspg-hexbinary'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oipf.dae.svg+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.dae.xhtml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.mippvcontrolmessage+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.pae.gem'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oipf.spdiscovery+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.spdlist+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.ueprofile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oipf.userprofile+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.olpc-sugar'] = MimeType{'iana',['xo'],false,''}
    data['application/vnd.oma-scws-config'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma-scws-http-request'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma-scws-http-response'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.bcast.associated-procedure-parameter+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.drm-trigger+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.imd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.ltkm'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.bcast.notification+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.provisioningtrigger'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.bcast.sgboot'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.bcast.sgdd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.sgdu'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.bcast.simple-symbol-container'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.bcast.smartcard-trigger+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.sprov+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.bcast.stkm'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.cab-address-book+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.cab-feature-handler+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.cab-pcc+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.cab-subs-invite+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.cab-user-prefs+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.dcd'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.dcdc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.dd2+xml'] = MimeType{'iana',['dd2'],true,''}
    data['application/vnd.oma.drm.risd+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.group-usage-list+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.lwm2m+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.lwm2m+tlv'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.pal+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.poc.detailed-progress-report+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.poc.final-report+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.poc.groups+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.poc.invocation-descriptor+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.poc.optimized-progress-report+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.push'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.oma.scidm.messages+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oma.xcap-directory+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.omads-email+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.omads-file+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.omads-folder+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.omaloc-supl-init'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.onepager'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.onepagertamp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.onepagertamx'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.onepagertat'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.onepagertatp'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.onepagertatx'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.openblox.game+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openblox.game-binary'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.openeye.oeb'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.openofficeorg.extension'] = MimeType{'apache',['oxt'],false,''}
    data['application/vnd.openstreetmap.data+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.custom-properties+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.customxmlproperties+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawing+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawingml.chart+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawingml.chartshapes+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawingml.diagramcolors+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawingml.diagramdata+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawingml.diagramlayout+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.drawingml.diagramstyle+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.extended-properties+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.commentauthors+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.comments+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.handoutmaster+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.notesmaster+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.notesslide+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.presentation'] = MimeType{'iana',['pptx'],false,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.presentation.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.presprops+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slide'] = MimeType{'iana',['sldx'],false,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slide+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slidelayout+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slidemaster+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slideshow'] = MimeType{'iana',['ppsx'],false,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slideshow.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.slideupdateinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.tablestyles+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.tags+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.template'] = MimeType{'iana',['potx'],false,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.template.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.presentationml.viewprops+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.calcchain+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.chartsheet+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.comments+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.connections+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.dialogsheet+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.externallink+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.pivotcachedefinition+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.pivotcacherecords+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.pivottable+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.querytable+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.revisionheaders+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.revisionlog+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.sharedstrings+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.sheet'] = MimeType{'iana',['xlsx'],false,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.sheet.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.sheetmetadata+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.styles+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.table+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.tablesinglecells+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.template'] = MimeType{'iana',['xltx'],false,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.template.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.usernames+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.volatiledependencies+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.spreadsheetml.worksheet+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.theme+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.themeoverride+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.vmldrawing'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.comments+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.document'] = MimeType{'iana',['docx'],false,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.document.glossary+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.document.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.endnotes+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.fonttable+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.footer+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.footnotes+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.numbering+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.settings+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.styles+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.template'] = MimeType{'iana',['dotx'],false,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.template.main+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-officedocument.wordprocessingml.websettings+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-package.core-properties+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-package.digital-signature-xmlsignature+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.openxmlformats-package.relationships+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oracle.resource+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.orange.indata'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.osa.netdeploy'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.osgeo.mapguide.package'] = MimeType{'iana',['mgp'],false,''}
    data['application/vnd.osgi.bundle'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.osgi.dp'] = MimeType{'iana',['dp'],false,''}
    data['application/vnd.osgi.subsystem'] = MimeType{'iana',['esa'],false,''}
    data['application/vnd.otps.ct-kip+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.oxli.countgraph'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.pagerduty+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.palm'] = MimeType{'iana',['pdb', 'pqa', 'oprc'],false,''}
    data['application/vnd.panoply'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.paos.xml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.patentdive'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.patientecommsdoc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.pawaafile'] = MimeType{'iana',['paw'],false,''}
    data['application/vnd.pcos'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.pg.format'] = MimeType{'iana',['str'],false,''}
    data['application/vnd.pg.osasli'] = MimeType{'iana',['ei6'],false,''}
    data['application/vnd.piaccess.application-licence'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.picsel'] = MimeType{'iana',['efif'],false,''}
    data['application/vnd.pmi.widget'] = MimeType{'iana',['wg'],false,''}
    data['application/vnd.poc.group-advertisement+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.pocketlearn'] = MimeType{'iana',['plf'],false,''}
    data['application/vnd.powerbuilder6'] = MimeType{'iana',['pbd'],false,''}
    data['application/vnd.powerbuilder6-s'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.powerbuilder7'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.powerbuilder7-s'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.powerbuilder75'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.powerbuilder75-s'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.preminet'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.previewsystems.box'] = MimeType{'iana',['box'],false,''}
    data['application/vnd.proteus.magazine'] = MimeType{'iana',['mgz'],false,''}
    data['application/vnd.psfs'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.publishare-delta-tree'] = MimeType{'iana',['qps'],false,''}
    data['application/vnd.pvi.ptid1'] = MimeType{'iana',['ptid'],false,''}
    data['application/vnd.pwg-multiplexed'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.pwg-xhtml-print+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.qualcomm.brew-app-res'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.quarantainenet'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.quark.quarkxpress'] = MimeType{'iana',['qxd', 'qxt', 'qwd', 'qwt', 'qxl', 'qxb'],false,''}
    data['application/vnd.quobject-quoxdocument'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.radisys.moml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-audit+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-audit-conf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-audit-conn+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-audit-dialog+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-audit-stream+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-conf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog-base+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog-fax-detect+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog-fax-sendrecv+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog-group+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog-speech+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.radisys.msml-dialog-transform+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.rainstor.data'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.rapid'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.rar'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.realvnc.bed'] = MimeType{'iana',['bed'],false,''}
    data['application/vnd.recordare.musicxml'] = MimeType{'iana',['mxl'],false,''}
    data['application/vnd.recordare.musicxml+xml'] = MimeType{'iana',['musicxml'],true,''}
    data['application/vnd.renlearn.rlprint'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.restful+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.rig.cryptonote'] = MimeType{'iana',['cryptonote'],false,''}
    data['application/vnd.rim.cod'] = MimeType{'apache',['cod'],false,''}
    data['application/vnd.rn-realmedia'] = MimeType{'apache',['rm'],false,''}
    data['application/vnd.rn-realmedia-vbr'] = MimeType{'apache',['rmvb'],false,''}
    data['application/vnd.route66.link66+xml'] = MimeType{'iana',['link66'],true,''}
    data['application/vnd.rs-274x'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ruckus.download'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.s3sms'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sailingtracker.track'] = MimeType{'iana',['st'],false,''}
    data['application/vnd.sbm.cid'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sbm.mid2'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.scribus'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.3df'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.csf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.doc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.eml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.mht'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.net'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.ppt'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.tiff'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealed.xls'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealedmedia.softseal.html'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sealedmedia.softseal.pdf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.seemail'] = MimeType{'iana',['see'],false,''}
    data['application/vnd.sema'] = MimeType{'iana',['sema'],false,''}
    data['application/vnd.semd'] = MimeType{'iana',['semd'],false,''}
    data['application/vnd.semf'] = MimeType{'iana',['semf'],false,''}
    data['application/vnd.shana.informed.formdata'] = MimeType{'iana',['ifm'],false,''}
    data['application/vnd.shana.informed.formtemplate'] = MimeType{'iana',['itp'],false,''}
    data['application/vnd.shana.informed.interchange'] = MimeType{'iana',['iif'],false,''}
    data['application/vnd.shana.informed.package'] = MimeType{'iana',['ipk'],false,''}
    data['application/vnd.shootproof+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.sigrok.session'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.simtech-mindmapper'] = MimeType{'iana',['twd', 'twds'],false,''}
    data['application/vnd.siren+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.smaf'] = MimeType{'iana',['mmf'],false,''}
    data['application/vnd.smart.notebook'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.smart.teacher'] = MimeType{'iana',['teacher'],false,''}
    data['application/vnd.software602.filler.form+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.software602.filler.form-xml-zip'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.solent.sdkm+xml'] = MimeType{'iana',['sdkm', 'sdkd'],true,''}
    data['application/vnd.spotfire.dxp'] = MimeType{'iana',['dxp'],false,''}
    data['application/vnd.spotfire.sfs'] = MimeType{'iana',['sfs'],false,''}
    data['application/vnd.sqlite3'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sss-cod'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sss-dtf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sss-ntf'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.stardivision.calc'] = MimeType{'apache',['sdc'],false,''}
    data['application/vnd.stardivision.draw'] = MimeType{'apache',['sda'],false,''}
    data['application/vnd.stardivision.impress'] = MimeType{'apache',['sdd'],false,''}
    data['application/vnd.stardivision.math'] = MimeType{'apache',['smf'],false,''}
    data['application/vnd.stardivision.writer'] = MimeType{'apache',['sdw', 'vor'],false,''}
    data['application/vnd.stardivision.writer-global'] = MimeType{'apache',['sgl'],false,''}
    data['application/vnd.stepmania.package'] = MimeType{'iana',['smzip'],false,''}
    data['application/vnd.stepmania.stepchart'] = MimeType{'iana',['sm'],false,''}
    data['application/vnd.street-stream'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.sun.wadl+xml'] = MimeType{'iana',['wadl'],true,''}
    data['application/vnd.sun.xml.calc'] = MimeType{'apache',['sxc'],false,''}
    data['application/vnd.sun.xml.calc.template'] = MimeType{'apache',['stc'],false,''}
    data['application/vnd.sun.xml.draw'] = MimeType{'apache',['sxd'],false,''}
    data['application/vnd.sun.xml.draw.template'] = MimeType{'apache',['std'],false,''}
    data['application/vnd.sun.xml.impress'] = MimeType{'apache',['sxi'],false,''}
    data['application/vnd.sun.xml.impress.template'] = MimeType{'apache',['sti'],false,''}
    data['application/vnd.sun.xml.math'] = MimeType{'apache',['sxm'],false,''}
    data['application/vnd.sun.xml.writer'] = MimeType{'apache',['sxw'],false,''}
    data['application/vnd.sun.xml.writer.global'] = MimeType{'apache',['sxg'],false,''}
    data['application/vnd.sun.xml.writer.template'] = MimeType{'apache',['stw'],false,''}
    data['application/vnd.sus-calendar'] = MimeType{'iana',['sus', 'susp'],false,''}
    data['application/vnd.svd'] = MimeType{'iana',['svd'],false,''}
    data['application/vnd.swiftview-ics'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.symbian.install'] = MimeType{'apache',['sis', 'sisx'],false,''}
    data['application/vnd.syncml+xml'] = MimeType{'iana',['xsm'],true,''}
    data['application/vnd.syncml.dm+wbxml'] = MimeType{'iana',['bdm'],false,''}
    data['application/vnd.syncml.dm+xml'] = MimeType{'iana',['xdm'],true,''}
    data['application/vnd.syncml.dm.notification'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.syncml.dmddf+wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.syncml.dmddf+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.syncml.dmtnds+wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.syncml.dmtnds+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.syncml.ds.notification'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.tableschema+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.tao.intent-module-archive'] = MimeType{'iana',['tao'],false,''}
    data['application/vnd.tcpdump.pcap'] = MimeType{'iana',['pcap', 'cap', 'dmp'],false,''}
    data['application/vnd.think-cell.ppttc+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.tmd.mediaflex.api+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.tml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.tmobile-livetv'] = MimeType{'iana',['tmo'],false,''}
    data['application/vnd.tri.onesource'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.trid.tpt'] = MimeType{'iana',['tpt'],false,''}
    data['application/vnd.triscape.mxs'] = MimeType{'iana',['mxs'],false,''}
    data['application/vnd.trueapp'] = MimeType{'iana',['tra'],false,''}
    data['application/vnd.truedoc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ubisoft.webplayer'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.ufdl'] = MimeType{'iana',['ufd', 'ufdl'],false,''}
    data['application/vnd.uiq.theme'] = MimeType{'iana',['utz'],false,''}
    data['application/vnd.umajin'] = MimeType{'iana',['umj'],false,''}
    data['application/vnd.unity'] = MimeType{'iana',['unityweb'],false,''}
    data['application/vnd.uoml+xml'] = MimeType{'iana',['uoml'],true,''}
    data['application/vnd.uplanet.alert'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.alert-wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.bearer-choice'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.bearer-choice-wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.cacheop'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.cacheop-wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.channel'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.channel-wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.list'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.list-wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.listcmd'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.listcmd-wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uplanet.signal'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.uri-map'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.valve.source.material'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.vcx'] = MimeType{'iana',['vcx'],false,''}
    data['application/vnd.vd-study'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.vectorworks'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.vel+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.verimatrix.vcas'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.veryant.thin'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.vidsoft.vidconference'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.visio'] = MimeType{'iana',['vsd', 'vst', 'vss', 'vsw'],false,''}
    data['application/vnd.visionary'] = MimeType{'iana',['vis'],false,''}
    data['application/vnd.vividence.scriptfile'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.vsf'] = MimeType{'iana',['vsf'],false,''}
    data['application/vnd.wap.sic'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wap.slc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wap.wbxml'] = MimeType{'iana',['wbxml'],false,''}
    data['application/vnd.wap.wmlc'] = MimeType{'iana',['wmlc'],false,''}
    data['application/vnd.wap.wmlscriptc'] = MimeType{'iana',['wmlsc'],false,''}
    data['application/vnd.webturbo'] = MimeType{'iana',['wtb'],false,''}
    data['application/vnd.wfa.p2p'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wfa.wsc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.windows.devicepairing'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wmc'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wmf.bootstrap'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wolfram.mathematica'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wolfram.mathematica.package'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wolfram.player'] = MimeType{'iana',['nbp'],false,''}
    data['application/vnd.wordperfect'] = MimeType{'iana',['wpd'],false,''}
    data['application/vnd.wqd'] = MimeType{'iana',['wqd'],false,''}
    data['application/vnd.wrq-hp3000-labelled'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wt.stf'] = MimeType{'iana',['stf'],false,''}
    data['application/vnd.wv.csp+wbxml'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.wv.csp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.wv.ssp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.xacml+json'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.xara'] = MimeType{'iana',['xar'],false,''}
    data['application/vnd.xfdl'] = MimeType{'iana',['xfdl'],false,''}
    data['application/vnd.xfdl.webform'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.xmi+xml'] = MimeType{'iana',[]string,true,''}
    data['application/vnd.xmpie.cpkg'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.xmpie.dpkg'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.xmpie.plan'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.xmpie.ppkg'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.xmpie.xlim'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.yamaha.hv-dic'] = MimeType{'iana',['hvd'],false,''}
    data['application/vnd.yamaha.hv-script'] = MimeType{'iana',['hvs'],false,''}
    data['application/vnd.yamaha.hv-voice'] = MimeType{'iana',['hvp'],false,''}
    data['application/vnd.yamaha.openscoreformat'] = MimeType{'iana',['osf'],false,''}
    data['application/vnd.yamaha.openscoreformat.osfpvg+xml'] = MimeType{'iana',['osfpvg'],true,''}
    data['application/vnd.yamaha.remote-setup'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.yamaha.smaf-audio'] = MimeType{'iana',['saf'],false,''}
    data['application/vnd.yamaha.smaf-phrase'] = MimeType{'iana',['spf'],false,''}
    data['application/vnd.yamaha.through-ngn'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.yamaha.tunnel-udpencap'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.yaoweme'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.yellowriver-custom-menu'] = MimeType{'iana',['cmp'],false,''}
    data['application/vnd.youtube.yt'] = MimeType{'iana',[]string,false,''}
    data['application/vnd.zul'] = MimeType{'iana',['zir', 'zirz'],false,''}
    data['application/vnd.zzazz.deck+xml'] = MimeType{'iana',['zaz'],true,''}
    data['application/voicexml+xml'] = MimeType{'iana',['vxml'],true,''}
    data['application/voucher-cms+json'] = MimeType{'iana',[]string,true,''}
    data['application/vq-rtcpxr'] = MimeType{'iana',[]string,false,''}
    data['application/wasm'] = MimeType{'',['wasm'],true,''}
    data['application/watcherinfo+xml'] = MimeType{'iana',[]string,true,''}
    data['application/webpush-options+json'] = MimeType{'iana',[]string,true,''}
    data['application/whoispp-query'] = MimeType{'iana',[]string,false,''}
    data['application/whoispp-response'] = MimeType{'iana',[]string,false,''}
    data['application/widget'] = MimeType{'iana',['wgt'],false,''}
    data['application/winhlp'] = MimeType{'apache',['hlp'],false,''}
    data['application/wita'] = MimeType{'iana',[]string,false,''}
    data['application/wordperfect5.1'] = MimeType{'iana',[]string,false,''}
    data['application/wsdl+xml'] = MimeType{'iana',['wsdl'],true,''}
    data['application/wspolicy+xml'] = MimeType{'iana',['wspolicy'],true,''}
    data['application/x-7z-compressed'] = MimeType{'apache',['7z'],false,''}
    data['application/x-abiword'] = MimeType{'apache',['abw'],false,''}
    data['application/x-ace-compressed'] = MimeType{'apache',['ace'],false,''}
    data['application/x-amf'] = MimeType{'apache',[]string,false,''}
    data['application/x-apple-diskimage'] = MimeType{'apache',['dmg'],false,''}
    data['application/x-arj'] = MimeType{'',['arj'],false,''}
    data['application/x-authorware-bin'] = MimeType{'apache',['aab', 'x32', 'u32', 'vox'],false,''}
    data['application/x-authorware-map'] = MimeType{'apache',['aam'],false,''}
    data['application/x-authorware-seg'] = MimeType{'apache',['aas'],false,''}
    data['application/x-bcpio'] = MimeType{'apache',['bcpio'],false,''}
    data['application/x-bdoc'] = MimeType{'',['bdoc'],false,''}
    data['application/x-bittorrent'] = MimeType{'apache',['torrent'],false,''}
    data['application/x-blorb'] = MimeType{'apache',['blb', 'blorb'],false,''}
    data['application/x-bzip'] = MimeType{'apache',['bz'],false,''}
    data['application/x-bzip2'] = MimeType{'apache',['bz2', 'boz'],false,''}
    data['application/x-cbr'] = MimeType{'apache',['cbr', 'cba', 'cbt', 'cbz', 'cb7'],false,''}
    data['application/x-cdlink'] = MimeType{'apache',['vcd'],false,''}
    data['application/x-cfs-compressed'] = MimeType{'apache',['cfs'],false,''}
    data['application/x-chat'] = MimeType{'apache',['chat'],false,''}
    data['application/x-chess-pgn'] = MimeType{'apache',['pgn'],false,''}
    data['application/x-chrome-extension'] = MimeType{'',['crx'],false,''}
    data['application/x-cocoa'] = MimeType{'nginx',['cco'],false,''}
    data['application/x-compress'] = MimeType{'apache',[]string,false,''}
    data['application/x-conference'] = MimeType{'apache',['nsc'],false,''}
    data['application/x-cpio'] = MimeType{'apache',['cpio'],false,''}
    data['application/x-csh'] = MimeType{'apache',['csh'],false,''}
    data['application/x-deb'] = MimeType{'',[]string,false,''}
    data['application/x-debian-package'] = MimeType{'apache',['deb', 'udeb'],false,''}
    data['application/x-dgc-compressed'] = MimeType{'apache',['dgc'],false,''}
    data['application/x-director'] = MimeType{'apache',['dir', 'dcr', 'dxr', 'cst', 'cct', 'cxt', 'w3d', 'fgd', 'swa'],false,''}
    data['application/x-doom'] = MimeType{'apache',['wad'],false,''}
    data['application/x-dtbncx+xml'] = MimeType{'apache',['ncx'],true,''}
    data['application/x-dtbook+xml'] = MimeType{'apache',['dtb'],true,''}
    data['application/x-dtbresource+xml'] = MimeType{'apache',['res'],true,''}
    data['application/x-dvi'] = MimeType{'apache',['dvi'],false,''}
    data['application/x-envoy'] = MimeType{'apache',['evy'],false,''}
    data['application/x-eva'] = MimeType{'apache',['eva'],false,''}
    data['application/x-font-bdf'] = MimeType{'apache',['bdf'],false,''}
    data['application/x-font-dos'] = MimeType{'apache',[]string,false,''}
    data['application/x-font-framemaker'] = MimeType{'apache',[]string,false,''}
    data['application/x-font-ghostscript'] = MimeType{'apache',['gsf'],false,''}
    data['application/x-font-libgrx'] = MimeType{'apache',[]string,false,''}
    data['application/x-font-linux-psf'] = MimeType{'apache',['psf'],false,''}
    data['application/x-font-pcf'] = MimeType{'apache',['pcf'],false,''}
    data['application/x-font-snf'] = MimeType{'apache',['snf'],false,''}
    data['application/x-font-speedo'] = MimeType{'apache',[]string,false,''}
    data['application/x-font-sunos-news'] = MimeType{'apache',[]string,false,''}
    data['application/x-font-type1'] = MimeType{'apache',['pfa', 'pfb', 'pfm', 'afm'],false,''}
    data['application/x-font-vfont'] = MimeType{'apache',[]string,false,''}
    data['application/x-freearc'] = MimeType{'apache',['arc'],false,''}
    data['application/x-futuresplash'] = MimeType{'apache',['spl'],false,''}
    data['application/x-gca-compressed'] = MimeType{'apache',['gca'],false,''}
    data['application/x-glulx'] = MimeType{'apache',['ulx'],false,''}
    data['application/x-gnumeric'] = MimeType{'apache',['gnumeric'],false,''}
    data['application/x-gramps-xml'] = MimeType{'apache',['gramps'],false,''}
    data['application/x-gtar'] = MimeType{'apache',['gtar'],false,''}
    data['application/x-gzip'] = MimeType{'apache',[]string,false,''}
    data['application/x-hdf'] = MimeType{'apache',['hdf'],false,''}
    data['application/x-httpd-php'] = MimeType{'',['php'],true,''}
    data['application/x-install-instructions'] = MimeType{'apache',['install'],false,''}
    data['application/x-iso9660-image'] = MimeType{'apache',['iso'],false,''}
    data['application/x-java-archive-diff'] = MimeType{'nginx',['jardiff'],false,''}
    data['application/x-java-jnlp-file'] = MimeType{'apache',['jnlp'],false,''}
    data['application/x-javascript'] = MimeType{'',[]string,true,''}
    data['application/x-latex'] = MimeType{'apache',['latex'],false,''}
    data['application/x-lua-bytecode'] = MimeType{'',['luac'],false,''}
    data['application/x-lzh-compressed'] = MimeType{'apache',['lzh', 'lha'],false,''}
    data['application/x-makeself'] = MimeType{'nginx',['run'],false,''}
    data['application/x-mie'] = MimeType{'apache',['mie'],false,''}
    data['application/x-mobipocket-ebook'] = MimeType{'apache',['prc', 'mobi'],false,''}
    data['application/x-mpegurl'] = MimeType{'',[]string,false,''}
    data['application/x-ms-application'] = MimeType{'apache',['application'],false,''}
    data['application/x-ms-shortcut'] = MimeType{'apache',['lnk'],false,''}
    data['application/x-ms-wmd'] = MimeType{'apache',['wmd'],false,''}
    data['application/x-ms-wmz'] = MimeType{'apache',['wmz'],false,''}
    data['application/x-ms-xbap'] = MimeType{'apache',['xbap'],false,''}
    data['application/x-msaccess'] = MimeType{'apache',['mdb'],false,''}
    data['application/x-msbinder'] = MimeType{'apache',['obd'],false,''}
    data['application/x-mscardfile'] = MimeType{'apache',['crd'],false,''}
    data['application/x-msclip'] = MimeType{'apache',['clp'],false,''}
    data['application/x-msdos-program'] = MimeType{'',['exe'],false,''}
    data['application/x-msdownload'] = MimeType{'apache',['exe', 'dll', 'com', 'bat', 'msi'],false,''}
    data['application/x-msmediaview'] = MimeType{'apache',['mvb', 'm13', 'm14'],false,''}
    data['application/x-msmetafile'] = MimeType{'apache',['wmf', 'wmz', 'emf', 'emz'],false,''}
    data['application/x-msmoney'] = MimeType{'apache',['mny'],false,''}
    data['application/x-mspublisher'] = MimeType{'apache',['pub'],false,''}
    data['application/x-msschedule'] = MimeType{'apache',['scd'],false,''}
    data['application/x-msterminal'] = MimeType{'apache',['trm'],false,''}
    data['application/x-mswrite'] = MimeType{'apache',['wri'],false,''}
    data['application/x-netcdf'] = MimeType{'apache',['nc', 'cdf'],false,''}
    data['application/x-ns-proxy-autoconfig'] = MimeType{'',['pac'],true,''}
    data['application/x-nzb'] = MimeType{'apache',['nzb'],false,''}
    data['application/x-perl'] = MimeType{'nginx',['pl', 'pm'],false,''}
    data['application/x-pilot'] = MimeType{'nginx',['prc', 'pdb'],false,''}
    data['application/x-pkcs12'] = MimeType{'apache',['p12', 'pfx'],false,''}
    data['application/x-pkcs7-certificates'] = MimeType{'apache',['p7b', 'spc'],false,''}
    data['application/x-pkcs7-certreqresp'] = MimeType{'apache',['p7r'],false,''}
    data['application/x-rar-compressed'] = MimeType{'apache',['rar'],false,''}
    data['application/x-redhat-package-manager'] = MimeType{'nginx',['rpm'],false,''}
    data['application/x-research-info-systems'] = MimeType{'apache',['ris'],false,''}
    data['application/x-sea'] = MimeType{'nginx',['sea'],false,''}
    data['application/x-sh'] = MimeType{'apache',['sh'],true,''}
    data['application/x-shar'] = MimeType{'apache',['shar'],false,''}
    data['application/x-shockwave-flash'] = MimeType{'apache',['swf'],false,''}
    data['application/x-silverlight-app'] = MimeType{'apache',['xap'],false,''}
    data['application/x-sql'] = MimeType{'apache',['sql'],false,''}
    data['application/x-stuffit'] = MimeType{'apache',['sit'],false,''}
    data['application/x-stuffitx'] = MimeType{'apache',['sitx'],false,''}
    data['application/x-subrip'] = MimeType{'apache',['srt'],false,''}
    data['application/x-sv4cpio'] = MimeType{'apache',['sv4cpio'],false,''}
    data['application/x-sv4crc'] = MimeType{'apache',['sv4crc'],false,''}
    data['application/x-t3vm-image'] = MimeType{'apache',['t3'],false,''}
    data['application/x-tads'] = MimeType{'apache',['gam'],false,''}
    data['application/x-tar'] = MimeType{'apache',['tar'],true,''}
    data['application/x-tcl'] = MimeType{'apache',['tcl', 'tk'],false,''}
    data['application/x-tex'] = MimeType{'apache',['tex'],false,''}
    data['application/x-tex-tfm'] = MimeType{'apache',['tfm'],false,''}
    data['application/x-texinfo'] = MimeType{'apache',['texinfo', 'texi'],false,''}
    data['application/x-tgif'] = MimeType{'apache',['obj'],false,''}
    data['application/x-ustar'] = MimeType{'apache',['ustar'],false,''}
    data['application/x-virtualbox-hdd'] = MimeType{'',['hdd'],true,''}
    data['application/x-virtualbox-ova'] = MimeType{'',['ova'],true,''}
    data['application/x-virtualbox-ovf'] = MimeType{'',['ovf'],true,''}
    data['application/x-virtualbox-vbox'] = MimeType{'',['vbox'],true,''}
    data['application/x-virtualbox-vbox-extpack'] = MimeType{'',['vbox-extpack'],false,''}
    data['application/x-virtualbox-vdi'] = MimeType{'',['vdi'],true,''}
    data['application/x-virtualbox-vhd'] = MimeType{'',['vhd'],true,''}
    data['application/x-virtualbox-vmdk'] = MimeType{'',['vmdk'],true,''}
    data['application/x-wais-source'] = MimeType{'apache',['src'],false,''}
    data['application/x-web-app-manifest+json'] = MimeType{'',['webapp'],true,''}
    data['application/x-www-form-urlencoded'] = MimeType{'iana',[]string,true,''}
    data['application/x-x509-ca-cert'] = MimeType{'apache',['der', 'crt', 'pem'],false,''}
    data['application/x-xfig'] = MimeType{'apache',['fig'],false,''}
    data['application/x-xliff+xml'] = MimeType{'apache',['xlf'],true,''}
    data['application/x-xpinstall'] = MimeType{'apache',['xpi'],false,''}
    data['application/x-xz'] = MimeType{'apache',['xz'],false,''}
    data['application/x-zmachine'] = MimeType{'apache',['z1', 'z2', 'z3', 'z4', 'z5', 'z6', 'z7', 'z8'],false,''}
    data['application/x400-bp'] = MimeType{'iana',[]string,false,''}
    data['application/xacml+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xaml+xml'] = MimeType{'apache',['xaml'],true,''}
    data['application/xcap-att+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xcap-caps+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xcap-diff+xml'] = MimeType{'iana',['xdf'],true,''}
    data['application/xcap-el+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xcap-error+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xcap-ns+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xcon-conference-info+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xcon-conference-info-diff+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xenc+xml'] = MimeType{'iana',['xenc'],true,''}
    data['application/xhtml+xml'] = MimeType{'iana',['xhtml', 'xht'],true,''}
    data['application/xhtml-voice+xml'] = MimeType{'apache',[]string,true,''}
    data['application/xliff+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xml'] = MimeType{'iana',['xml', 'xsl', 'xsd', 'rng'],true,''}
    data['application/xml-dtd'] = MimeType{'iana',['dtd'],true,''}
    data['application/xml-external-parsed-entity'] = MimeType{'iana',[]string,false,''}
    data['application/xml-patch+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xmpp+xml'] = MimeType{'iana',[]string,true,''}
    data['application/xop+xml'] = MimeType{'iana',['xop'],true,''}
    data['application/xproc+xml'] = MimeType{'apache',['xpl'],true,''}
    data['application/xslt+xml'] = MimeType{'iana',['xslt'],true,''}
    data['application/xspf+xml'] = MimeType{'apache',['xspf'],true,''}
    data['application/xv+xml'] = MimeType{'iana',['mxml', 'xhvml', 'xvml', 'xvm'],true,''}
    data['application/yang'] = MimeType{'iana',['yang'],false,''}
    data['application/yang-data+json'] = MimeType{'iana',[]string,true,''}
    data['application/yang-data+xml'] = MimeType{'iana',[]string,true,''}
    data['application/yang-patch+json'] = MimeType{'iana',[]string,true,''}
    data['application/yang-patch+xml'] = MimeType{'iana',[]string,true,''}
    data['application/yin+xml'] = MimeType{'iana',['yin'],true,''}
    data['application/zip'] = MimeType{'iana',['zip'],false,''}
    data['application/zlib'] = MimeType{'iana',[]string,false,''}
    data['application/zstd'] = MimeType{'iana',[]string,false,''}
    data['audio/1d-interleaved-parityfec'] = MimeType{'iana',[]string,false,''}
    data['audio/32kadpcm'] = MimeType{'iana',[]string,false,''}
    data['audio/3gpp'] = MimeType{'iana',['3gpp'],false,''}
    data['audio/3gpp2'] = MimeType{'iana',[]string,false,''}
    data['audio/aac'] = MimeType{'iana',[]string,false,''}
    data['audio/ac3'] = MimeType{'iana',[]string,false,''}
    data['audio/adpcm'] = MimeType{'apache',['adp'],false,''}
    data['audio/amr'] = MimeType{'iana',[]string,false,''}
    data['audio/amr-wb'] = MimeType{'iana',[]string,false,''}
    data['audio/amr-wb+'] = MimeType{'iana',[]string,false,''}
    data['audio/aptx'] = MimeType{'iana',[]string,false,''}
    data['audio/asc'] = MimeType{'iana',[]string,false,''}
    data['audio/atrac-advanced-lossless'] = MimeType{'iana',[]string,false,''}
    data['audio/atrac-x'] = MimeType{'iana',[]string,false,''}
    data['audio/atrac3'] = MimeType{'iana',[]string,false,''}
    data['audio/basic'] = MimeType{'iana',['au', 'snd'],false,''}
    data['audio/bv16'] = MimeType{'iana',[]string,false,''}
    data['audio/bv32'] = MimeType{'iana',[]string,false,''}
    data['audio/clearmode'] = MimeType{'iana',[]string,false,''}
    data['audio/cn'] = MimeType{'iana',[]string,false,''}
    data['audio/dat12'] = MimeType{'iana',[]string,false,''}
    data['audio/dls'] = MimeType{'iana',[]string,false,''}
    data['audio/dsr-es201108'] = MimeType{'iana',[]string,false,''}
    data['audio/dsr-es202050'] = MimeType{'iana',[]string,false,''}
    data['audio/dsr-es202211'] = MimeType{'iana',[]string,false,''}
    data['audio/dsr-es202212'] = MimeType{'iana',[]string,false,''}
    data['audio/dv'] = MimeType{'iana',[]string,false,''}
    data['audio/dvi4'] = MimeType{'iana',[]string,false,''}
    data['audio/eac3'] = MimeType{'iana',[]string,false,''}
    data['audio/encaprtp'] = MimeType{'iana',[]string,false,''}
    data['audio/evrc'] = MimeType{'iana',[]string,false,''}
    data['audio/evrc-qcp'] = MimeType{'iana',[]string,false,''}
    data['audio/evrc0'] = MimeType{'iana',[]string,false,''}
    data['audio/evrc1'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcb'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcb0'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcb1'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcnw'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcnw0'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcnw1'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcwb'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcwb0'] = MimeType{'iana',[]string,false,''}
    data['audio/evrcwb1'] = MimeType{'iana',[]string,false,''}
    data['audio/evs'] = MimeType{'iana',[]string,false,''}
    data['audio/fwdred'] = MimeType{'iana',[]string,false,''}
    data['audio/g711-0'] = MimeType{'iana',[]string,false,''}
    data['audio/g719'] = MimeType{'iana',[]string,false,''}
    data['audio/g722'] = MimeType{'iana',[]string,false,''}
    data['audio/g7221'] = MimeType{'iana',[]string,false,''}
    data['audio/g723'] = MimeType{'iana',[]string,false,''}
    data['audio/g726-16'] = MimeType{'iana',[]string,false,''}
    data['audio/g726-24'] = MimeType{'iana',[]string,false,''}
    data['audio/g726-32'] = MimeType{'iana',[]string,false,''}
    data['audio/g726-40'] = MimeType{'iana',[]string,false,''}
    data['audio/g728'] = MimeType{'iana',[]string,false,''}
    data['audio/g729'] = MimeType{'iana',[]string,false,''}
    data['audio/g7291'] = MimeType{'iana',[]string,false,''}
    data['audio/g729d'] = MimeType{'iana',[]string,false,''}
    data['audio/g729e'] = MimeType{'iana',[]string,false,''}
    data['audio/gsm'] = MimeType{'iana',[]string,false,''}
    data['audio/gsm-efr'] = MimeType{'iana',[]string,false,''}
    data['audio/gsm-hr-08'] = MimeType{'iana',[]string,false,''}
    data['audio/ilbc'] = MimeType{'iana',[]string,false,''}
    data['audio/ip-mr_v2.5'] = MimeType{'iana',[]string,false,''}
    data['audio/isac'] = MimeType{'apache',[]string,false,''}
    data['audio/l16'] = MimeType{'iana',[]string,false,''}
    data['audio/l20'] = MimeType{'iana',[]string,false,''}
    data['audio/l24'] = MimeType{'iana',[]string,false,''}
    data['audio/l8'] = MimeType{'iana',[]string,false,''}
    data['audio/lpc'] = MimeType{'iana',[]string,false,''}
    data['audio/melp'] = MimeType{'iana',[]string,false,''}
    data['audio/melp1200'] = MimeType{'iana',[]string,false,''}
    data['audio/melp2400'] = MimeType{'iana',[]string,false,''}
    data['audio/melp600'] = MimeType{'iana',[]string,false,''}
    data['audio/midi'] = MimeType{'apache',['mid', 'midi', 'kar', 'rmi'],false,''}
    data['audio/mobile-xmf'] = MimeType{'iana',[]string,false,''}
    data['audio/mp3'] = MimeType{'',['mp3'],false,''}
    data['audio/mp4'] = MimeType{'iana',['m4a', 'mp4a'],false,''}
    data['audio/mp4a-latm'] = MimeType{'iana',[]string,false,''}
    data['audio/mpa'] = MimeType{'iana',[]string,false,''}
    data['audio/mpa-robust'] = MimeType{'iana',[]string,false,''}
    data['audio/mpeg'] = MimeType{'iana',['mpga', 'mp2', 'mp2a', 'mp3', 'm2a', 'm3a'],false,''}
    data['audio/mpeg4-generic'] = MimeType{'iana',[]string,false,''}
    data['audio/musepack'] = MimeType{'apache',[]string,false,''}
    data['audio/ogg'] = MimeType{'iana',['oga', 'ogg', 'spx'],false,''}
    data['audio/opus'] = MimeType{'iana',[]string,false,''}
    data['audio/parityfec'] = MimeType{'iana',[]string,false,''}
    data['audio/pcma'] = MimeType{'iana',[]string,false,''}
    data['audio/pcma-wb'] = MimeType{'iana',[]string,false,''}
    data['audio/pcmu'] = MimeType{'iana',[]string,false,''}
    data['audio/pcmu-wb'] = MimeType{'iana',[]string,false,''}
    data['audio/prs.sid'] = MimeType{'iana',[]string,false,''}
    data['audio/qcelp'] = MimeType{'iana',[]string,false,''}
    data['audio/raptorfec'] = MimeType{'iana',[]string,false,''}
    data['audio/red'] = MimeType{'iana',[]string,false,''}
    data['audio/rtp-enc-aescm128'] = MimeType{'iana',[]string,false,''}
    data['audio/rtp-midi'] = MimeType{'iana',[]string,false,''}
    data['audio/rtploopback'] = MimeType{'iana',[]string,false,''}
    data['audio/rtx'] = MimeType{'iana',[]string,false,''}
    data['audio/s3m'] = MimeType{'apache',['s3m'],false,''}
    data['audio/silk'] = MimeType{'apache',['sil'],false,''}
    data['audio/smv'] = MimeType{'iana',[]string,false,''}
    data['audio/smv-qcp'] = MimeType{'iana',[]string,false,''}
    data['audio/smv0'] = MimeType{'iana',[]string,false,''}
    data['audio/sp-midi'] = MimeType{'iana',[]string,false,''}
    data['audio/speex'] = MimeType{'iana',[]string,false,''}
    data['audio/t140c'] = MimeType{'iana',[]string,false,''}
    data['audio/t38'] = MimeType{'iana',[]string,false,''}
    data['audio/telephone-event'] = MimeType{'iana',[]string,false,''}
    data['audio/tetra_acelp'] = MimeType{'iana',[]string,false,''}
    data['audio/tone'] = MimeType{'iana',[]string,false,''}
    data['audio/uemclip'] = MimeType{'iana',[]string,false,''}
    data['audio/ulpfec'] = MimeType{'iana',[]string,false,''}
    data['audio/usac'] = MimeType{'iana',[]string,false,''}
    data['audio/vdvi'] = MimeType{'iana',[]string,false,''}
    data['audio/vmr-wb'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.3gpp.iufp'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.4sb'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.audiokoz'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.celp'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.cisco.nse'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.cmles.radio-events'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.cns.anp1'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.cns.inf1'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dece.audio'] = MimeType{'iana',['uva', 'uvva'],false,''}
    data['audio/vnd.digital-winds'] = MimeType{'iana',['eol'],false,''}
    data['audio/vnd.dlna.adts'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.heaac.1'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.heaac.2'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.mlp'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.mps'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.pl2'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.pl2x'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.pl2z'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dolby.pulse.1'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dra'] = MimeType{'iana',['dra'],false,''}
    data['audio/vnd.dts'] = MimeType{'iana',['dts'],false,''}
    data['audio/vnd.dts.hd'] = MimeType{'iana',['dtshd'],false,''}
    data['audio/vnd.dts.uhd'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.dvb.file'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.everad.plj'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.hns.audio'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.lucent.voice'] = MimeType{'iana',['lvp'],false,''}
    data['audio/vnd.ms-playready.media.pya'] = MimeType{'iana',['pya'],false,''}
    data['audio/vnd.nokia.mobile-xmf'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.nortel.vbk'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.nuera.ecelp4800'] = MimeType{'iana',['ecelp4800'],false,''}
    data['audio/vnd.nuera.ecelp7470'] = MimeType{'iana',['ecelp7470'],false,''}
    data['audio/vnd.nuera.ecelp9600'] = MimeType{'iana',['ecelp9600'],false,''}
    data['audio/vnd.octel.sbc'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.presonus.multitrack'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.qcelp'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.rhetorex.32kadpcm'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.rip'] = MimeType{'iana',['rip'],false,''}
    data['audio/vnd.rn-realaudio'] = MimeType{'',[]string,false,''}
    data['audio/vnd.sealedmedia.softseal.mpeg'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.vmx.cvsd'] = MimeType{'iana',[]string,false,''}
    data['audio/vnd.wave'] = MimeType{'',[]string,false,''}
    data['audio/vorbis'] = MimeType{'iana',[]string,false,''}
    data['audio/vorbis-config'] = MimeType{'iana',[]string,false,''}
    data['audio/wav'] = MimeType{'',['wav'],false,''}
    data['audio/wave'] = MimeType{'',['wav'],false,''}
    data['audio/webm'] = MimeType{'apache',['weba'],false,''}
    data['audio/x-aac'] = MimeType{'apache',['aac'],false,''}
    data['audio/x-aiff'] = MimeType{'apache',['aif', 'aiff', 'aifc'],false,''}
    data['audio/x-caf'] = MimeType{'apache',['caf'],false,''}
    data['audio/x-flac'] = MimeType{'apache',['flac'],false,''}
    data['audio/x-m4a'] = MimeType{'nginx',['m4a'],false,''}
    data['audio/x-matroska'] = MimeType{'apache',['mka'],false,''}
    data['audio/x-mpegurl'] = MimeType{'apache',['m3u'],false,''}
    data['audio/x-ms-wax'] = MimeType{'apache',['wax'],false,''}
    data['audio/x-ms-wma'] = MimeType{'apache',['wma'],false,''}
    data['audio/x-pn-realaudio'] = MimeType{'apache',['ram', 'ra'],false,''}
    data['audio/x-pn-realaudio-plugin'] = MimeType{'apache',['rmp'],false,''}
    data['audio/x-realaudio'] = MimeType{'nginx',['ra'],false,''}
    data['audio/x-tta'] = MimeType{'apache',[]string,false,''}
    data['audio/x-wav'] = MimeType{'apache',['wav'],false,''}
    data['audio/xm'] = MimeType{'apache',['xm'],false,''}
    data['chemical/x-cdx'] = MimeType{'apache',['cdx'],false,''}
    data['chemical/x-cif'] = MimeType{'apache',['cif'],false,''}
    data['chemical/x-cmdf'] = MimeType{'apache',['cmdf'],false,''}
    data['chemical/x-cml'] = MimeType{'apache',['cml'],false,''}
    data['chemical/x-csml'] = MimeType{'apache',['csml'],false,''}
    data['chemical/x-pdb'] = MimeType{'apache',[]string,false,''}
    data['chemical/x-xyz'] = MimeType{'apache',['xyz'],false,''}
    data['font/collection'] = MimeType{'iana',['ttc'],false,''}
    data['font/otf'] = MimeType{'iana',['otf'],true,''}
    data['font/sfnt'] = MimeType{'iana',[]string,false,''}
    data['font/ttf'] = MimeType{'iana',['ttf'],false,''}
    data['font/woff'] = MimeType{'iana',['woff'],false,''}
    data['font/woff2'] = MimeType{'iana',['woff2'],false,''}
    data['image/aces'] = MimeType{'iana',['exr'],false,''}
    data['image/apng'] = MimeType{'',['apng'],false,''}
    data['image/avci'] = MimeType{'iana',[]string,false,''}
    data['image/avcs'] = MimeType{'iana',[]string,false,''}
    data['image/bmp'] = MimeType{'iana',['bmp'],true,''}
    data['image/cgm'] = MimeType{'iana',['cgm'],false,''}
    data['image/dicom-rle'] = MimeType{'iana',['drle'],false,''}
    data['image/emf'] = MimeType{'iana',['emf'],false,''}
    data['image/fits'] = MimeType{'iana',['fits'],false,''}
    data['image/g3fax'] = MimeType{'iana',['g3'],false,''}
    data['image/gif'] = MimeType{'iana',['gif'],false,''}
    data['image/heic'] = MimeType{'iana',['heic'],false,''}
    data['image/heic-sequence'] = MimeType{'iana',['heics'],false,''}
    data['image/heif'] = MimeType{'iana',['heif'],false,''}
    data['image/heif-sequence'] = MimeType{'iana',['heifs'],false,''}
    data['image/ief'] = MimeType{'iana',['ief'],false,''}
    data['image/jls'] = MimeType{'iana',['jls'],false,''}
    data['image/jp2'] = MimeType{'iana',['jp2', 'jpg2'],false,''}
    data['image/jpeg'] = MimeType{'iana',['jpeg', 'jpg', 'jpe'],false,''}
    data['image/jpm'] = MimeType{'iana',['jpm'],false,''}
    data['image/jpx'] = MimeType{'iana',['jpx', 'jpf'],false,''}
    data['image/jxr'] = MimeType{'iana',['jxr'],false,''}
    data['image/ktx'] = MimeType{'iana',['ktx'],false,''}
    data['image/naplps'] = MimeType{'iana',[]string,false,''}
    data['image/pjpeg'] = MimeType{'',[]string,false,''}
    data['image/png'] = MimeType{'iana',['png'],false,''}
    data['image/prs.btif'] = MimeType{'iana',['btif'],false,''}
    data['image/prs.pti'] = MimeType{'iana',['pti'],false,''}
    data['image/pwg-raster'] = MimeType{'iana',[]string,false,''}
    data['image/sgi'] = MimeType{'apache',['sgi'],false,''}
    data['image/svg+xml'] = MimeType{'iana',['svg', 'svgz'],true,''}
    data['image/t38'] = MimeType{'iana',['t38'],false,''}
    data['image/tiff'] = MimeType{'iana',['tif', 'tiff'],false,''}
    data['image/tiff-fx'] = MimeType{'iana',['tfx'],false,''}
    data['image/vnd.adobe.photoshop'] = MimeType{'iana',['psd'],true,''}
    data['image/vnd.airzip.accelerator.azv'] = MimeType{'iana',['azv'],false,''}
    data['image/vnd.cns.inf2'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.dece.graphic'] = MimeType{'iana',['uvi', 'uvvi', 'uvg', 'uvvg'],false,''}
    data['image/vnd.djvu'] = MimeType{'iana',['djvu', 'djv'],false,''}
    data['image/vnd.dvb.subtitle'] = MimeType{'iana',['sub'],false,''}
    data['image/vnd.dwg'] = MimeType{'iana',['dwg'],false,''}
    data['image/vnd.dxf'] = MimeType{'iana',['dxf'],false,''}
    data['image/vnd.fastbidsheet'] = MimeType{'iana',['fbs'],false,''}
    data['image/vnd.fpx'] = MimeType{'iana',['fpx'],false,''}
    data['image/vnd.fst'] = MimeType{'iana',['fst'],false,''}
    data['image/vnd.fujixerox.edmics-mmr'] = MimeType{'iana',['mmr'],false,''}
    data['image/vnd.fujixerox.edmics-rlc'] = MimeType{'iana',['rlc'],false,''}
    data['image/vnd.globalgraphics.pgb'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.microsoft.icon'] = MimeType{'iana',['ico'],false,''}
    data['image/vnd.mix'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.mozilla.apng'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.ms-modi'] = MimeType{'iana',['mdi'],false,''}
    data['image/vnd.ms-photo'] = MimeType{'apache',['wdp'],false,''}
    data['image/vnd.net-fpx'] = MimeType{'iana',['npx'],false,''}
    data['image/vnd.radiance'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.sealed.png'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.sealedmedia.softseal.gif'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.sealedmedia.softseal.jpg'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.svf'] = MimeType{'iana',[]string,false,''}
    data['image/vnd.tencent.tap'] = MimeType{'iana',['tap'],false,''}
    data['image/vnd.valve.source.texture'] = MimeType{'iana',['vtf'],false,''}
    data['image/vnd.wap.wbmp'] = MimeType{'iana',['wbmp'],false,''}
    data['image/vnd.xiff'] = MimeType{'iana',['xif'],false,''}
    data['image/vnd.zbrush.pcx'] = MimeType{'iana',['pcx'],false,''}
    data['image/webp'] = MimeType{'apache',['webp'],false,''}
    data['image/wmf'] = MimeType{'iana',['wmf'],false,''}
    data['image/x-3ds'] = MimeType{'apache',['3ds'],false,''}
    data['image/x-cmu-raster'] = MimeType{'apache',['ras'],false,''}
    data['image/x-cmx'] = MimeType{'apache',['cmx'],false,''}
    data['image/x-freehand'] = MimeType{'apache',['fh', 'fhc', 'fh4', 'fh5', 'fh7'],false,''}
    data['image/x-icon'] = MimeType{'apache',['ico'],true,''}
    data['image/x-jng'] = MimeType{'nginx',['jng'],false,''}
    data['image/x-mrsid-image'] = MimeType{'apache',['sid'],false,''}
    data['image/x-ms-bmp'] = MimeType{'nginx',['bmp'],true,''}
    data['image/x-pcx'] = MimeType{'apache',['pcx'],false,''}
    data['image/x-pict'] = MimeType{'apache',['pic', 'pct'],false,''}
    data['image/x-portable-anymap'] = MimeType{'apache',['pnm'],false,''}
    data['image/x-portable-bitmap'] = MimeType{'apache',['pbm'],false,''}
    data['image/x-portable-graymap'] = MimeType{'apache',['pgm'],false,''}
    data['image/x-portable-pixmap'] = MimeType{'apache',['ppm'],false,''}
    data['image/x-rgb'] = MimeType{'apache',['rgb'],false,''}
    data['image/x-tga'] = MimeType{'apache',['tga'],false,''}
    data['image/x-xbitmap'] = MimeType{'apache',['xbm'],false,''}
    data['image/x-xcf'] = MimeType{'',[]string,false,''}
    data['image/x-xpixmap'] = MimeType{'apache',['xpm'],false,''}
    data['image/x-xwindowdump'] = MimeType{'apache',['xwd'],false,''}
    data['message/cpim'] = MimeType{'iana',[]string,false,''}
    data['message/delivery-status'] = MimeType{'iana',[]string,false,''}
    data['message/disposition-notification'] = MimeType{'iana',['disposition-notification'],false,''}
    data['message/external-body'] = MimeType{'iana',[]string,false,''}
    data['message/feedback-report'] = MimeType{'iana',[]string,false,''}
    data['message/global'] = MimeType{'iana',['u8msg'],false,''}
    data['message/global-delivery-status'] = MimeType{'iana',['u8dsn'],false,''}
    data['message/global-disposition-notification'] = MimeType{'iana',['u8mdn'],false,''}
    data['message/global-headers'] = MimeType{'iana',['u8hdr'],false,''}
    data['message/http'] = MimeType{'iana',[]string,false,''}
    data['message/imdn+xml'] = MimeType{'iana',[]string,true,''}
    data['message/news'] = MimeType{'iana',[]string,false,''}
    data['message/partial'] = MimeType{'iana',[]string,false,''}
    data['message/rfc822'] = MimeType{'iana',['eml', 'mime'],true,''}
    data['message/s-http'] = MimeType{'iana',[]string,false,''}
    data['message/sip'] = MimeType{'iana',[]string,false,''}
    data['message/sipfrag'] = MimeType{'iana',[]string,false,''}
    data['message/tracking-status'] = MimeType{'iana',[]string,false,''}
    data['message/vnd.si.simp'] = MimeType{'iana',[]string,false,''}
    data['message/vnd.wfa.wsc'] = MimeType{'iana',['wsc'],false,''}
    data['model/3mf'] = MimeType{'iana',['3mf'],false,''}
    data['model/gltf+json'] = MimeType{'iana',['gltf'],true,''}
    data['model/gltf-binary'] = MimeType{'iana',['glb'],true,''}
    data['model/iges'] = MimeType{'iana',['igs', 'iges'],false,''}
    data['model/mesh'] = MimeType{'iana',['msh', 'mesh', 'silo'],false,''}
    data['model/stl'] = MimeType{'iana',['stl'],false,''}
    data['model/vnd.collada+xml'] = MimeType{'iana',['dae'],true,''}
    data['model/vnd.dwf'] = MimeType{'iana',['dwf'],false,''}
    data['model/vnd.flatland.3dml'] = MimeType{'iana',[]string,false,''}
    data['model/vnd.gdl'] = MimeType{'iana',['gdl'],false,''}
    data['model/vnd.gs-gdl'] = MimeType{'apache',[]string,false,''}
    data['model/vnd.gs.gdl'] = MimeType{'iana',[]string,false,''}
    data['model/vnd.gtw'] = MimeType{'iana',['gtw'],false,''}
    data['model/vnd.moml+xml'] = MimeType{'iana',[]string,true,''}
    data['model/vnd.mts'] = MimeType{'iana',['mts'],false,''}
    data['model/vnd.opengex'] = MimeType{'iana',['ogex'],false,''}
    data['model/vnd.parasolid.transmit.binary'] = MimeType{'iana',['x_b'],false,''}
    data['model/vnd.parasolid.transmit.text'] = MimeType{'iana',['x_t'],false,''}
    data['model/vnd.rosette.annotated-data-model'] = MimeType{'iana',[]string,false,''}
    data['model/vnd.usdz+zip'] = MimeType{'iana',['usdz'],false,''}
    data['model/vnd.valve.source.compiled-map'] = MimeType{'iana',['bsp'],false,''}
    data['model/vnd.vtu'] = MimeType{'iana',['vtu'],false,''}
    data['model/vrml'] = MimeType{'iana',['wrl', 'vrml'],false,''}
    data['model/x3d+binary'] = MimeType{'apache',['x3db', 'x3dbz'],false,''}
    data['model/x3d+fastinfoset'] = MimeType{'iana',['x3db'],false,''}
    data['model/x3d+vrml'] = MimeType{'apache',['x3dv', 'x3dvz'],false,''}
    data['model/x3d+xml'] = MimeType{'iana',['x3d', 'x3dz'],true,''}
    data['model/x3d-vrml'] = MimeType{'iana',['x3dv'],false,''}
    data['multipart/alternative'] = MimeType{'iana',[]string,false,''}
    data['multipart/appledouble'] = MimeType{'iana',[]string,false,''}
    data['multipart/byteranges'] = MimeType{'iana',[]string,false,''}
    data['multipart/digest'] = MimeType{'iana',[]string,false,''}
    data['multipart/encrypted'] = MimeType{'iana',[]string,false,''}
    data['multipart/form-data'] = MimeType{'iana',[]string,false,''}
    data['multipart/header-set'] = MimeType{'iana',[]string,false,''}
    data['multipart/mixed'] = MimeType{'iana',[]string,false,''}
    data['multipart/multilingual'] = MimeType{'iana',[]string,false,''}
    data['multipart/parallel'] = MimeType{'iana',[]string,false,''}
    data['multipart/related'] = MimeType{'iana',[]string,false,''}
    data['multipart/report'] = MimeType{'iana',[]string,false,''}
    data['multipart/signed'] = MimeType{'iana',[]string,false,''}
    data['multipart/vnd.bint.med-plus'] = MimeType{'iana',[]string,false,''}
    data['multipart/voice-message'] = MimeType{'iana',[]string,false,''}
    data['multipart/x-mixed-replace'] = MimeType{'iana',[]string,false,''}
    data['text/1d-interleaved-parityfec'] = MimeType{'iana',[]string,false,''}
    data['text/cache-manifest'] = MimeType{'iana',['appcache', 'manifest'],true,''}
    data['text/calendar'] = MimeType{'iana',['ics', 'ifb'],false,''}
    data['text/calender'] = MimeType{'',[]string,true,''}
    data['text/cmd'] = MimeType{'',[]string,true,''}
    data['text/coffeescript'] = MimeType{'',['coffee', 'litcoffee'],false,''}
    data['text/css'] = MimeType{'iana',['css'],true,'UTF-8'}
    data['text/csv'] = MimeType{'iana',['csv'],true,''}
    data['text/csv-schema'] = MimeType{'iana',[]string,false,''}
    data['text/directory'] = MimeType{'iana',[]string,false,''}
    data['text/dns'] = MimeType{'iana',[]string,false,''}
    data['text/ecmascript'] = MimeType{'iana',[]string,false,''}
    data['text/encaprtp'] = MimeType{'iana',[]string,false,''}
    data['text/enriched'] = MimeType{'iana',[]string,false,''}
    data['text/fwdred'] = MimeType{'iana',[]string,false,''}
    data['text/grammar-ref-list'] = MimeType{'iana',[]string,false,''}
    data['text/html'] = MimeType{'iana',['html', 'htm', 'shtml'],true,''}
    data['text/jade'] = MimeType{'',['jade'],false,''}
    data['text/javascript'] = MimeType{'iana',[]string,true,''}
    data['text/jcr-cnd'] = MimeType{'iana',[]string,false,''}
    data['text/jsx'] = MimeType{'',['jsx'],true,''}
    data['text/less'] = MimeType{'',['less'],true,''}
    data['text/markdown'] = MimeType{'iana',['markdown', 'md'],true,''}
    data['text/mathml'] = MimeType{'nginx',['mml'],false,''}
    data['text/mdx'] = MimeType{'',['mdx'],true,''}
    data['text/mizar'] = MimeType{'iana',[]string,false,''}
    data['text/n3'] = MimeType{'iana',['n3'],true,''}
    data['text/parameters'] = MimeType{'iana',[]string,false,''}
    data['text/parityfec'] = MimeType{'iana',[]string,false,''}
    data['text/plain'] = MimeType{'iana',['txt', 'text', 'conf', 'def', 'list', 'log', 'in', 'ini'],true,''}
    data['text/provenance-notation'] = MimeType{'iana',[]string,false,''}
    data['text/prs.fallenstein.rst'] = MimeType{'iana',[]string,false,''}
    data['text/prs.lines.tag'] = MimeType{'iana',['dsc'],false,''}
    data['text/prs.prop.logic'] = MimeType{'iana',[]string,false,''}
    data['text/raptorfec'] = MimeType{'iana',[]string,false,''}
    data['text/red'] = MimeType{'iana',[]string,false,''}
    data['text/rfc822-headers'] = MimeType{'iana',[]string,false,''}
    data['text/richtext'] = MimeType{'iana',['rtx'],true,''}
    data['text/rtf'] = MimeType{'iana',['rtf'],true,''}
    data['text/rtp-enc-aescm128'] = MimeType{'iana',[]string,false,''}
    data['text/rtploopback'] = MimeType{'iana',[]string,false,''}
    data['text/rtx'] = MimeType{'iana',[]string,false,''}
    data['text/sgml'] = MimeType{'iana',['sgml', 'sgm'],false,''}
    data['text/shex'] = MimeType{'',['shex'],false,''}
    data['text/slim'] = MimeType{'',['slim', 'slm'],false,''}
    data['text/strings'] = MimeType{'iana',[]string,false,''}
    data['text/stylus'] = MimeType{'',['stylus', 'styl'],false,''}
    data['text/t140'] = MimeType{'iana',[]string,false,''}
    data['text/tab-separated-values'] = MimeType{'iana',['tsv'],true,''}
    data['text/troff'] = MimeType{'iana',['t', 'tr', 'roff', 'man', 'me', 'ms'],false,''}
    data['text/turtle'] = MimeType{'iana',['ttl'],false,'UTF-8'}
    data['text/ulpfec'] = MimeType{'iana',[]string,false,''}
    data['text/uri-list'] = MimeType{'iana',['uri', 'uris', 'urls'],true,''}
    data['text/vcard'] = MimeType{'iana',['vcard'],true,''}
    data['text/vnd.a'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.abc'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.ascii-art'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.curl'] = MimeType{'iana',['curl'],false,''}
    data['text/vnd.curl.dcurl'] = MimeType{'apache',['dcurl'],false,''}
    data['text/vnd.curl.mcurl'] = MimeType{'apache',['mcurl'],false,''}
    data['text/vnd.curl.scurl'] = MimeType{'apache',['scurl'],false,''}
    data['text/vnd.debian.copyright'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.dmclientscript'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.dvb.subtitle'] = MimeType{'iana',['sub'],false,''}
    data['text/vnd.esmertec.theme-descriptor'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.fly'] = MimeType{'iana',['fly'],false,''}
    data['text/vnd.fmi.flexstor'] = MimeType{'iana',['flx'],false,''}
    data['text/vnd.gml'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.graphviz'] = MimeType{'iana',['gv'],false,''}
    data['text/vnd.hgl'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.in3d.3dml'] = MimeType{'iana',['3dml'],false,''}
    data['text/vnd.in3d.spot'] = MimeType{'iana',['spot'],false,''}
    data['text/vnd.iptc.newsml'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.iptc.nitf'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.latex-z'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.motorola.reflex'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.ms-mediapackage'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.net2phone.commcenter.command'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.radisys.msml-basic-layout'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.senx.warpscript'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.si.uricatalogue'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.sun.j2me.app-descriptor'] = MimeType{'iana',['jad'],false,''}
    data['text/vnd.trolltech.linguist'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.wap.si'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.wap.sl'] = MimeType{'iana',[]string,false,''}
    data['text/vnd.wap.wml'] = MimeType{'iana',['wml'],false,''}
    data['text/vnd.wap.wmlscript'] = MimeType{'iana',['wmls'],false,''}
    data['text/vtt'] = MimeType{'',['vtt'],true,'UTF-8'}
    data['text/x-asm'] = MimeType{'apache',['s', 'asm'],false,''}
    data['text/x-c'] = MimeType{'apache',['c', 'cc', 'cxx', 'cpp', 'h', 'hh', 'dic'],false,''}
    data['text/x-component'] = MimeType{'nginx',['htc'],false,''}
    data['text/x-fortran'] = MimeType{'apache',['f', 'for', 'f77', 'f90'],false,''}
    data['text/x-gwt-rpc'] = MimeType{'',[]string,true,''}
    data['text/x-handlebars-template'] = MimeType{'',['hbs'],false,''}
    data['text/x-java-source'] = MimeType{'apache',['java'],false,''}
    data['text/x-jquery-tmpl'] = MimeType{'',[]string,true,''}
    data['text/x-lua'] = MimeType{'',['lua'],false,''}
    data['text/x-markdown'] = MimeType{'',['mkd'],true,''}
    data['text/x-nfo'] = MimeType{'apache',['nfo'],false,''}
    data['text/x-opml'] = MimeType{'apache',['opml'],false,''}
    data['text/x-org'] = MimeType{'',['org'],true,''}
    data['text/x-pascal'] = MimeType{'apache',['p', 'pas'],false,''}
    data['text/x-processing'] = MimeType{'',['pde'],true,''}
    data['text/x-sass'] = MimeType{'',['sass'],false,''}
    data['text/x-scss'] = MimeType{'',['scss'],false,''}
    data['text/x-setext'] = MimeType{'apache',['etx'],false,''}
    data['text/x-sfv'] = MimeType{'apache',['sfv'],false,''}
    data['text/x-suse-ymp'] = MimeType{'',['ymp'],true,''}
    data['text/x-uuencode'] = MimeType{'apache',['uu'],false,''}
    data['text/x-vcalendar'] = MimeType{'apache',['vcs'],false,''}
    data['text/x-vcard'] = MimeType{'apache',['vcf'],false,''}
    data['text/xml'] = MimeType{'iana',['xml'],true,''}
    data['text/xml-external-parsed-entity'] = MimeType{'iana',[]string,false,''}
    data['text/yaml'] = MimeType{'',['yaml', 'yml'],false,''}
    data['video/1d-interleaved-parityfec'] = MimeType{'iana',[]string,false,''}
    data['video/3gpp'] = MimeType{'iana',['3gp', '3gpp'],false,''}
    data['video/3gpp-tt'] = MimeType{'iana',[]string,false,''}
    data['video/3gpp2'] = MimeType{'iana',['3g2'],false,''}
    data['video/bmpeg'] = MimeType{'iana',[]string,false,''}
    data['video/bt656'] = MimeType{'iana',[]string,false,''}
    data['video/celb'] = MimeType{'iana',[]string,false,''}
    data['video/dv'] = MimeType{'iana',[]string,false,''}
    data['video/encaprtp'] = MimeType{'iana',[]string,false,''}
    data['video/h261'] = MimeType{'iana',['h261'],false,''}
    data['video/h263'] = MimeType{'iana',['h263'],false,''}
    data['video/h263-1998'] = MimeType{'iana',[]string,false,''}
    data['video/h263-2000'] = MimeType{'iana',[]string,false,''}
    data['video/h264'] = MimeType{'iana',['h264'],false,''}
    data['video/h264-rcdo'] = MimeType{'iana',[]string,false,''}
    data['video/h264-svc'] = MimeType{'iana',[]string,false,''}
    data['video/h265'] = MimeType{'iana',[]string,false,''}
    data['video/iso.segment'] = MimeType{'iana',[]string,false,''}
    data['video/jpeg'] = MimeType{'iana',['jpgv'],false,''}
    data['video/jpeg2000'] = MimeType{'iana',[]string,false,''}
    data['video/jpm'] = MimeType{'apache',['jpm', 'jpgm'],false,''}
    data['video/mj2'] = MimeType{'iana',['mj2', 'mjp2'],false,''}
    data['video/mp1s'] = MimeType{'iana',[]string,false,''}
    data['video/mp2p'] = MimeType{'iana',[]string,false,''}
    data['video/mp2t'] = MimeType{'iana',['ts'],false,''}
    data['video/mp4'] = MimeType{'iana',['mp4', 'mp4v', 'mpg4'],false,''}
    data['video/mp4v-es'] = MimeType{'iana',[]string,false,''}
    data['video/mpeg'] = MimeType{'iana',['mpeg', 'mpg', 'mpe', 'm1v', 'm2v'],false,''}
    data['video/mpeg4-generic'] = MimeType{'iana',[]string,false,''}
    data['video/mpv'] = MimeType{'iana',[]string,false,''}
    data['video/nv'] = MimeType{'iana',[]string,false,''}
    data['video/ogg'] = MimeType{'iana',['ogv'],false,''}
    data['video/parityfec'] = MimeType{'iana',[]string,false,''}
    data['video/pointer'] = MimeType{'iana',[]string,false,''}
    data['video/quicktime'] = MimeType{'iana',['qt', 'mov'],false,''}
    data['video/raptorfec'] = MimeType{'iana',[]string,false,''}
    data['video/raw'] = MimeType{'iana',[]string,false,''}
    data['video/rtp-enc-aescm128'] = MimeType{'iana',[]string,false,''}
    data['video/rtploopback'] = MimeType{'iana',[]string,false,''}
    data['video/rtx'] = MimeType{'iana',[]string,false,''}
    data['video/smpte291'] = MimeType{'iana',[]string,false,''}
    data['video/smpte292m'] = MimeType{'iana',[]string,false,''}
    data['video/ulpfec'] = MimeType{'iana',[]string,false,''}
    data['video/vc1'] = MimeType{'iana',[]string,false,''}
    data['video/vc2'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.cctv'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.dece.hd'] = MimeType{'iana',['uvh', 'uvvh'],false,''}
    data['video/vnd.dece.mobile'] = MimeType{'iana',['uvm', 'uvvm'],false,''}
    data['video/vnd.dece.mp4'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.dece.pd'] = MimeType{'iana',['uvp', 'uvvp'],false,''}
    data['video/vnd.dece.sd'] = MimeType{'iana',['uvs', 'uvvs'],false,''}
    data['video/vnd.dece.video'] = MimeType{'iana',['uvv', 'uvvv'],false,''}
    data['video/vnd.directv.mpeg'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.directv.mpeg-tts'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.dlna.mpeg-tts'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.dvb.file'] = MimeType{'iana',['dvb'],false,''}
    data['video/vnd.fvt'] = MimeType{'iana',['fvt'],false,''}
    data['video/vnd.hns.video'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.iptvforum.1dparityfec-1010'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.iptvforum.1dparityfec-2005'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.iptvforum.2dparityfec-1010'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.iptvforum.2dparityfec-2005'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.iptvforum.ttsavc'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.iptvforum.ttsmpeg2'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.motorola.video'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.motorola.videop'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.mpegurl'] = MimeType{'iana',['mxu', 'm4u'],false,''}
    data['video/vnd.ms-playready.media.pyv'] = MimeType{'iana',['pyv'],false,''}
    data['video/vnd.nokia.interleaved-multimedia'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.nokia.mp4vr'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.nokia.videovoip'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.objectvideo'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.radgamettools.bink'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.radgamettools.smacker'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.sealed.mpeg1'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.sealed.mpeg4'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.sealed.swf'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.sealedmedia.softseal.mov'] = MimeType{'iana',[]string,false,''}
    data['video/vnd.uvvu.mp4'] = MimeType{'iana',['uvu', 'uvvu'],false,''}
    data['video/vnd.vivo'] = MimeType{'iana',['viv'],false,''}
    data['video/vp8'] = MimeType{'iana',[]string,false,''}
    data['video/webm'] = MimeType{'apache',['webm'],false,''}
    data['video/x-f4v'] = MimeType{'apache',['f4v'],false,''}
    data['video/x-fli'] = MimeType{'apache',['fli'],false,''}
    data['video/x-flv'] = MimeType{'apache',['flv'],false,''}
    data['video/x-m4v'] = MimeType{'apache',['m4v'],false,''}
    data['video/x-matroska'] = MimeType{'apache',['mkv', 'mk3d', 'mks'],false,''}
    data['video/x-mng'] = MimeType{'apache',['mng'],false,''}
    data['video/x-ms-asf'] = MimeType{'apache',['asf', 'asx'],false,''}
    data['video/x-ms-vob'] = MimeType{'apache',['vob'],false,''}
    data['video/x-ms-wm'] = MimeType{'apache',['wm'],false,''}
    data['video/x-ms-wmv'] = MimeType{'apache',['wmv'],false,''}
    data['video/x-ms-wmx'] = MimeType{'apache',['wmx'],false,''}
    data['video/x-ms-wvx'] = MimeType{'apache',['wvx'],false,''}
    data['video/x-msvideo'] = MimeType{'apache',['avi'],false,''}
    data['video/x-sgi-movie'] = MimeType{'apache',['movie'],false,''}
    data['video/x-smv'] = MimeType{'apache',['smv'],false,''}
    data['x-conference/x-cooltalk'] = MimeType{'apache',['ice'],false,''}
    data['x-shader/x-fragment'] = MimeType{'',[]string,true,''}
    data['x-shader/x-vertex'] = MimeType{'',[]string,true,''}
    return data
}